// Copyright (C) 1991-2013 Altera Corporation
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, Altera MegaCore Function License 
// Agreement, or other applicable license agreement, including, 
// without limitation, that your use is for the sole purpose of 
// programming logic devices manufactured by Altera and sold by 
// Altera or its authorized distributors.  Please refer to the 
// applicable agreement for further details.

// VENDOR "Altera"
// PROGRAM "Quartus II 64-Bit"
// VERSION "Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Full Version"

// DATE "12/09/2016 18:33:53"

// 
// Device: Altera EP4CE115F29C8 Package FBGA780
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module system (
	altera_reserved_tms,
	altera_reserved_tck,
	altera_reserved_tdi,
	altera_reserved_tdo,
	CLK,
	nRST,
	\syif.halt ,
	\syif.load ,
	\syif.addr ,
	\syif.store ,
	\syif.REN ,
	\syif.WEN ,
	\syif.tbCTRL );
input 	altera_reserved_tms;
input 	altera_reserved_tck;
input 	altera_reserved_tdi;
output 	altera_reserved_tdo;
input 	CLK;
input 	nRST;
output 	\syif.halt ;
output 	[31:0] \syif.load ;
input 	[31:0] \syif.addr ;
input 	[31:0] \syif.store ;
input 	\syif.REN ;
input 	\syif.WEN ;
input 	\syif.tbCTRL ;

// Design Ports Information
// syif.halt	=>  Location: PIN_AC10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[0]	=>  Location: PIN_AC11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[1]	=>  Location: PIN_AD12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[2]	=>  Location: PIN_AB13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[3]	=>  Location: PIN_AB10,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[4]	=>  Location: PIN_AB2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[5]	=>  Location: PIN_AE18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[6]	=>  Location: PIN_V1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[7]	=>  Location: PIN_AD14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[8]	=>  Location: PIN_AG22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[9]	=>  Location: PIN_U28,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[10]	=>  Location: PIN_D14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[11]	=>  Location: PIN_AD15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[12]	=>  Location: PIN_J15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[13]	=>  Location: PIN_C14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[14]	=>  Location: PIN_Y14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[15]	=>  Location: PIN_R5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[16]	=>  Location: PIN_AB15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[17]	=>  Location: PIN_B17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[18]	=>  Location: PIN_C13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[19]	=>  Location: PIN_D13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[20]	=>  Location: PIN_A12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[21]	=>  Location: PIN_AF16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[22]	=>  Location: PIN_D16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[23]	=>  Location: PIN_AH17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[24]	=>  Location: PIN_AC15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[25]	=>  Location: PIN_V2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[26]	=>  Location: PIN_AB1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[27]	=>  Location: PIN_Y15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[28]	=>  Location: PIN_AH23,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[29]	=>  Location: PIN_AC14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[30]	=>  Location: PIN_AF18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.load[31]	=>  Location: PIN_T25,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[1]	=>  Location: PIN_AG15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.tbCTRL	=>  Location: PIN_AH15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[0]	=>  Location: PIN_AH18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[3]	=>  Location: PIN_AH19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[2]	=>  Location: PIN_H15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[5]	=>  Location: PIN_AC17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[4]	=>  Location: PIN_AG21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[7]	=>  Location: PIN_AG12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[6]	=>  Location: PIN_AH12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[9]	=>  Location: PIN_C12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[8]	=>  Location: PIN_AB16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[11]	=>  Location: PIN_AF15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[10]	=>  Location: PIN_AE15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[13]	=>  Location: PIN_J14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[12]	=>  Location: PIN_AA16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[15]	=>  Location: PIN_AA15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[14]	=>  Location: PIN_AG17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[23]	=>  Location: PIN_C15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[22]	=>  Location: PIN_AE17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.WEN	=>  Location: PIN_AD17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.REN	=>  Location: PIN_W22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[21]	=>  Location: PIN_C16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[29]	=>  Location: PIN_AE16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[28]	=>  Location: PIN_D15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[31]	=>  Location: PIN_F15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[30]	=>  Location: PIN_U21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[20]	=>  Location: PIN_AH21,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[17]	=>  Location: PIN_AG18,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[16]	=>  Location: PIN_U27,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[19]	=>  Location: PIN_AB14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[18]	=>  Location: PIN_V4,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[25]	=>  Location: PIN_AH22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[24]	=>  Location: PIN_AG19,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[27]	=>  Location: PIN_AF17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.addr[26]	=>  Location: PIN_A17,	 I/O Standard: 2.5 V,	 Current Strength: Default
// nRST	=>  Location: PIN_Y2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// CLK	=>  Location: PIN_J1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[0]	=>  Location: PIN_AF12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[1]	=>  Location: PIN_G14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[2]	=>  Location: PIN_Y12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[3]	=>  Location: PIN_Y13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[4]	=>  Location: PIN_AE13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[5]	=>  Location: PIN_W2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[6]	=>  Location: PIN_AE12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[7]	=>  Location: PIN_AB12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[8]	=>  Location: PIN_AC12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[9]	=>  Location: PIN_V3,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[10]	=>  Location: PIN_AF13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[11]	=>  Location: PIN_AA13,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[12]	=>  Location: PIN_D12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[13]	=>  Location: PIN_AA12,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[14]	=>  Location: PIN_H14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[15]	=>  Location: PIN_U2,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[16]	=>  Location: PIN_T7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[17]	=>  Location: PIN_AH11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[18]	=>  Location: PIN_E14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[19]	=>  Location: PIN_AE11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[20]	=>  Location: PIN_AF14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[21]	=>  Location: PIN_AE14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[22]	=>  Location: PIN_Y22,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[23]	=>  Location: PIN_AA14,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[24]	=>  Location: PIN_G15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[25]	=>  Location: PIN_U1,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[26]	=>  Location: PIN_AD11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[27]	=>  Location: PIN_E15,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[28]	=>  Location: PIN_H16,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[29]	=>  Location: PIN_AF11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[30]	=>  Location: PIN_U24,	 I/O Standard: 2.5 V,	 Current Strength: Default
// syif.store[31]	=>  Location: PIN_AG11,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tms	=>  Location: PIN_P8,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tck	=>  Location: PIN_P5,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdi	=>  Location: PIN_P7,	 I/O Standard: 2.5 V,	 Current Strength: Default
// altera_reserved_tdo	=>  Location: PIN_P6,	 I/O Standard: 2.5 V,	 Current Strength: Default


wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire \CPU|DP|prif.dmemren~q ;
wire \CPU|DP|prif.dmemwen~q ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ;
wire \RAM|LessThan1~0_combout ;
wire \ramaddr~0_combout ;
wire \ramaddr~1_combout ;
wire \ramaddr~2_combout ;
wire \ramaddr~3_combout ;
wire \ramaddr~4_combout ;
wire \ramaddr~5_combout ;
wire \ramaddr~6_combout ;
wire \ramaddr~7_combout ;
wire \ramaddr~8_combout ;
wire \ramaddr~9_combout ;
wire \ramaddr~10_combout ;
wire \ramaddr~11_combout ;
wire \ramaddr~12_combout ;
wire \ramaddr~13_combout ;
wire \ramaddr~14_combout ;
wire \ramaddr~15_combout ;
wire \ramaddr~16_combout ;
wire \ramaddr~17_combout ;
wire \ramaddr~18_combout ;
wire \ramaddr~19_combout ;
wire \ramaddr~20_combout ;
wire \ramaddr~21_combout ;
wire \ramaddr~22_combout ;
wire \ramaddr~23_combout ;
wire \ramaddr~24_combout ;
wire \ramaddr~25_combout ;
wire \ramaddr~26_combout ;
wire \ramaddr~27_combout ;
wire \ramaddr~28_combout ;
wire \ramaddr~29_combout ;
wire \ramaddr~30_combout ;
wire \ramaddr~31_combout ;
wire \ramaddr~32_combout ;
wire \ramaddr~33_combout ;
wire \ramaddr~34_combout ;
wire \ramaddr~35_combout ;
wire \ramWEN~0_combout ;
wire \ramREN~0_combout ;
wire \ramaddr~36_combout ;
wire \ramaddr~37_combout ;
wire \ramaddr~38_combout ;
wire \ramaddr~39_combout ;
wire \ramaddr~40_combout ;
wire \ramaddr~41_combout ;
wire \ramaddr~42_combout ;
wire \ramaddr~43_combout ;
wire \ramaddr~44_combout ;
wire \ramaddr~45_combout ;
wire \ramaddr~46_combout ;
wire \ramaddr~47_combout ;
wire \ramaddr~48_combout ;
wire \ramaddr~49_combout ;
wire \ramaddr~50_combout ;
wire \ramaddr~51_combout ;
wire \ramaddr~52_combout ;
wire \ramaddr~53_combout ;
wire \ramaddr~54_combout ;
wire \ramaddr~55_combout ;
wire \ramaddr~56_combout ;
wire \ramaddr~57_combout ;
wire \ramaddr~58_combout ;
wire \ramaddr~59_combout ;
wire \ramaddr~60_combout ;
wire \ramaddr~61_combout ;
wire \ramaddr~62_combout ;
wire \ramaddr~63_combout ;
wire \RAM|always0~21_combout ;
wire \RAM|always1~0_combout ;
wire \RAM|ramif.ramload[0]~0_combout ;
wire \RAM|ramif.ramload[1]~1_combout ;
wire \RAM|ramif.ramload[2]~2_combout ;
wire \RAM|ramif.ramload[3]~3_combout ;
wire \RAM|ramif.ramload[4]~4_combout ;
wire \RAM|ramif.ramload[5]~5_combout ;
wire \RAM|ramif.ramload[6]~6_combout ;
wire \RAM|ramif.ramload[7]~7_combout ;
wire \RAM|ramif.ramload[8]~8_combout ;
wire \RAM|ramif.ramload[9]~9_combout ;
wire \RAM|ramif.ramload[10]~10_combout ;
wire \RAM|ramif.ramload[11]~11_combout ;
wire \RAM|ramif.ramload[12]~12_combout ;
wire \RAM|ramif.ramload[13]~13_combout ;
wire \RAM|ramif.ramload[14]~14_combout ;
wire \RAM|ramif.ramload[15]~15_combout ;
wire \RAM|ramif.ramload[16]~16_combout ;
wire \RAM|ramif.ramload[17]~17_combout ;
wire \RAM|ramif.ramload[18]~18_combout ;
wire \RAM|ramif.ramload[19]~19_combout ;
wire \RAM|ramif.ramload[20]~20_combout ;
wire \RAM|ramif.ramload[21]~21_combout ;
wire \RAM|ramif.ramload[22]~22_combout ;
wire \RAM|ramif.ramload[23]~23_combout ;
wire \RAM|ramif.ramload[24]~24_combout ;
wire \RAM|ramif.ramload[25]~25_combout ;
wire \RAM|ramif.ramload[26]~26_combout ;
wire \RAM|ramif.ramload[27]~27_combout ;
wire \RAM|ramif.ramload[28]~28_combout ;
wire \RAM|ramif.ramload[29]~29_combout ;
wire \RAM|ramif.ramload[30]~30_combout ;
wire \RAM|ramif.ramload[31]~31_combout ;
wire \RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ;
wire \CPUCLK~q ;
wire \ramstore~0_combout ;
wire \ramstore~1_combout ;
wire \ramstore~2_combout ;
wire \ramstore~3_combout ;
wire \ramstore~4_combout ;
wire \ramstore~5_combout ;
wire \ramstore~6_combout ;
wire \ramstore~7_combout ;
wire \ramstore~8_combout ;
wire \ramstore~9_combout ;
wire \ramstore~10_combout ;
wire \ramstore~11_combout ;
wire \ramstore~12_combout ;
wire \ramstore~13_combout ;
wire \ramstore~14_combout ;
wire \ramstore~15_combout ;
wire \ramstore~16_combout ;
wire \ramstore~17_combout ;
wire \ramstore~18_combout ;
wire \ramstore~19_combout ;
wire \ramstore~20_combout ;
wire \ramstore~21_combout ;
wire \ramstore~22_combout ;
wire \ramstore~23_combout ;
wire \ramstore~24_combout ;
wire \ramstore~25_combout ;
wire \ramstore~26_combout ;
wire \ramstore~27_combout ;
wire \ramstore~28_combout ;
wire \ramstore~29_combout ;
wire \ramstore~30_combout ;
wire \ramstore~31_combout ;
wire \Equal0~0_combout ;
wire \CPUCLK~0_combout ;
wire \count[3]~0_combout ;
wire \count[2]~1_combout ;
wire \count[1]~2_combout ;
wire \count~3_combout ;
wire \ramaddr~29_wirecell_combout ;
wire \altera_internal_jtag~TCKUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~10 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ;
wire \auto_hub|~GND~combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ;
wire \syif.addr[1]~input_o ;
wire \syif.tbCTRL~input_o ;
wire \syif.addr[0]~input_o ;
wire \syif.addr[3]~input_o ;
wire \syif.addr[2]~input_o ;
wire \syif.addr[5]~input_o ;
wire \syif.addr[4]~input_o ;
wire \syif.addr[7]~input_o ;
wire \syif.addr[6]~input_o ;
wire \syif.addr[9]~input_o ;
wire \syif.addr[8]~input_o ;
wire \syif.addr[11]~input_o ;
wire \syif.addr[10]~input_o ;
wire \syif.addr[13]~input_o ;
wire \syif.addr[12]~input_o ;
wire \syif.addr[15]~input_o ;
wire \syif.addr[14]~input_o ;
wire \syif.addr[23]~input_o ;
wire \syif.addr[22]~input_o ;
wire \syif.WEN~input_o ;
wire \syif.REN~input_o ;
wire \syif.addr[21]~input_o ;
wire \syif.addr[29]~input_o ;
wire \syif.addr[28]~input_o ;
wire \syif.addr[31]~input_o ;
wire \syif.addr[30]~input_o ;
wire \syif.addr[20]~input_o ;
wire \syif.addr[17]~input_o ;
wire \syif.addr[16]~input_o ;
wire \syif.addr[19]~input_o ;
wire \syif.addr[18]~input_o ;
wire \syif.addr[25]~input_o ;
wire \syif.addr[24]~input_o ;
wire \syif.addr[27]~input_o ;
wire \syif.addr[26]~input_o ;
wire \nRST~input_o ;
wire \CLK~input_o ;
wire \syif.store[0]~input_o ;
wire \syif.store[1]~input_o ;
wire \syif.store[2]~input_o ;
wire \syif.store[3]~input_o ;
wire \syif.store[4]~input_o ;
wire \syif.store[5]~input_o ;
wire \syif.store[6]~input_o ;
wire \syif.store[7]~input_o ;
wire \syif.store[8]~input_o ;
wire \syif.store[9]~input_o ;
wire \syif.store[10]~input_o ;
wire \syif.store[11]~input_o ;
wire \syif.store[12]~input_o ;
wire \syif.store[13]~input_o ;
wire \syif.store[14]~input_o ;
wire \syif.store[15]~input_o ;
wire \syif.store[16]~input_o ;
wire \syif.store[17]~input_o ;
wire \syif.store[18]~input_o ;
wire \syif.store[19]~input_o ;
wire \syif.store[20]~input_o ;
wire \syif.store[21]~input_o ;
wire \syif.store[22]~input_o ;
wire \syif.store[23]~input_o ;
wire \syif.store[24]~input_o ;
wire \syif.store[25]~input_o ;
wire \syif.store[26]~input_o ;
wire \syif.store[27]~input_o ;
wire \syif.store[28]~input_o ;
wire \syif.store[29]~input_o ;
wire \syif.store[30]~input_o ;
wire \syif.store[31]~input_o ;
wire \altera_internal_jtag~TCKUTAPclkctrl_outclk ;
wire \CPUCLK~clkctrl_outclk ;
wire \nRST~inputclkctrl_outclk ;
wire \CLK~inputclkctrl_outclk ;
wire \CPU|DP|dpif.halt~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ;
wire \altera_reserved_tms~input_o ;
wire \altera_reserved_tck~input_o ;
wire \altera_reserved_tdi~input_o ;
wire \altera_internal_jtag~TDIUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ;
wire \altera_internal_jtag~TMSUTAP ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ;
wire \~QIC_CREATED_GND~I_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ;
wire \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ;
wire \altera_internal_jtag~TDO ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg ;
wire [9:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg ;
wire [5:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg ;
wire [2:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt ;
wire [15:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state ;
wire [4:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter ;
wire [3:0] \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR ;
wire [3:0] count;
wire [31:0] \CPU|DP|prif.dmemstore ;
wire [31:0] \CPU|DP|prif.dmemaddr ;
wire [31:0] \CPU|DP|pc ;
wire [3:0] \RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg ;


ram RAM(
	.is_in_use_reg(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.LessThan1(\RAM|LessThan1~0_combout ),
	.\ramif.ramaddr ({\ramaddr~43_combout ,\ramaddr~45_combout ,\ramaddr~39_combout ,\ramaddr~41_combout ,\ramaddr~61_combout ,\ramaddr~63_combout ,\ramaddr~57_combout ,gnd,\ramaddr~33_combout ,\ramaddr~35_combout ,\ramaddr~37_combout ,\ramaddr~47_combout ,\ramaddr~53_combout ,gnd,
\ramaddr~49_combout ,\ramaddr~51_combout ,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,gnd,\ramaddr~1_combout ,gnd}),
	.ramaddr(\ramaddr~3_combout ),
	.ramaddr1(\ramaddr~5_combout ),
	.ramaddr2(\ramaddr~7_combout ),
	.ramaddr3(\ramaddr~9_combout ),
	.ramaddr4(\ramaddr~11_combout ),
	.ramaddr5(\ramaddr~13_combout ),
	.ramaddr6(\ramaddr~15_combout ),
	.ramaddr7(\ramaddr~17_combout ),
	.ramaddr8(\ramaddr~19_combout ),
	.ramaddr9(\ramaddr~21_combout ),
	.ramaddr10(\ramaddr~23_combout ),
	.ramaddr11(\ramaddr~25_combout ),
	.ramaddr12(\ramaddr~27_combout ),
	.ramaddr13(\ramaddr~29_combout ),
	.ramaddr14(\ramaddr~31_combout ),
	.\ramif.ramWEN (\ramWEN~0_combout ),
	.\ramif.ramREN (\ramREN~0_combout ),
	.ramaddr15(\ramaddr~55_combout ),
	.ramaddr16(\ramaddr~59_combout ),
	.always0(\RAM|always0~21_combout ),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.ir_loaded_address_reg_0(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.ir_loaded_address_reg_1(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.ir_loaded_address_reg_2(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.ir_loaded_address_reg_3(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.tdo(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.ramstore(\ramstore~0_combout ),
	.ramstore1(\ramstore~1_combout ),
	.ramstore2(\ramstore~2_combout ),
	.ramstore3(\ramstore~3_combout ),
	.ramstore4(\ramstore~4_combout ),
	.ramstore5(\ramstore~5_combout ),
	.ramstore6(\ramstore~6_combout ),
	.ramstore7(\ramstore~7_combout ),
	.ramstore8(\ramstore~8_combout ),
	.ramstore9(\ramstore~9_combout ),
	.ramstore10(\ramstore~10_combout ),
	.ramstore11(\ramstore~11_combout ),
	.ramstore12(\ramstore~12_combout ),
	.ramstore13(\ramstore~13_combout ),
	.ramstore14(\ramstore~14_combout ),
	.ramstore15(\ramstore~15_combout ),
	.ramstore16(\ramstore~16_combout ),
	.ramstore17(\ramstore~17_combout ),
	.ramstore18(\ramstore~18_combout ),
	.ramstore19(\ramstore~19_combout ),
	.ramstore20(\ramstore~20_combout ),
	.ramstore21(\ramstore~21_combout ),
	.ramstore22(\ramstore~22_combout ),
	.ramstore23(\ramstore~23_combout ),
	.ramstore24(\ramstore~24_combout ),
	.ramstore25(\ramstore~25_combout ),
	.ramstore26(\ramstore~26_combout ),
	.ramstore27(\ramstore~27_combout ),
	.ramstore28(\ramstore~28_combout ),
	.ramstore29(\ramstore~29_combout ),
	.ramstore30(\ramstore~30_combout ),
	.ramstore31(\ramstore~31_combout ),
	.ramaddr17(\ramaddr~29_wirecell_combout ),
	.altera_internal_jtag(\altera_internal_jtag~TDIUTAP ),
	.state_4(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.irf_reg_0_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.irf_reg_1_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.irf_reg_2_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.irf_reg_3_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.irf_reg_4_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.node_ena_1(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.clr_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.virtual_ir_scan_reg(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.state_3(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.state_5(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.state_8(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.nRST(\nRST~input_o ),
	.altera_internal_jtag1(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.CLK(\CLK~inputclkctrl_outclk ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline CPU(
	.prifdmemaddr_1(\CPU|DP|prif.dmemaddr [1]),
	.pc_1(\CPU|DP|pc [1]),
	.prifdmemren(\CPU|DP|prif.dmemren~q ),
	.prifdmemwen(\CPU|DP|prif.dmemwen~q ),
	.prifdmemaddr_0(\CPU|DP|prif.dmemaddr [0]),
	.pc_0(\CPU|DP|pc [0]),
	.prifdmemaddr_3(\CPU|DP|prif.dmemaddr [3]),
	.prifdmemaddr_2(\CPU|DP|prif.dmemaddr [2]),
	.prifdmemaddr_5(\CPU|DP|prif.dmemaddr [5]),
	.prifdmemaddr_4(\CPU|DP|prif.dmemaddr [4]),
	.prifdmemaddr_7(\CPU|DP|prif.dmemaddr [7]),
	.prifdmemaddr_6(\CPU|DP|prif.dmemaddr [6]),
	.prifdmemaddr_9(\CPU|DP|prif.dmemaddr [9]),
	.prifdmemaddr_8(\CPU|DP|prif.dmemaddr [8]),
	.prifdmemaddr_11(\CPU|DP|prif.dmemaddr [11]),
	.prifdmemaddr_10(\CPU|DP|prif.dmemaddr [10]),
	.prifdmemaddr_13(\CPU|DP|prif.dmemaddr [13]),
	.prifdmemaddr_12(\CPU|DP|prif.dmemaddr [12]),
	.prifdmemaddr_15(\CPU|DP|prif.dmemaddr [15]),
	.prifdmemaddr_14(\CPU|DP|prif.dmemaddr [14]),
	.prifdmemaddr_23(\CPU|DP|prif.dmemaddr [23]),
	.prifdmemaddr_22(\CPU|DP|prif.dmemaddr [22]),
	.prifdmemaddr_21(\CPU|DP|prif.dmemaddr [21]),
	.prifdmemaddr_29(\CPU|DP|prif.dmemaddr [29]),
	.prifdmemaddr_28(\CPU|DP|prif.dmemaddr [28]),
	.prifdmemaddr_31(\CPU|DP|prif.dmemaddr [31]),
	.prifdmemaddr_30(\CPU|DP|prif.dmemaddr [30]),
	.prifdmemaddr_20(\CPU|DP|prif.dmemaddr [20]),
	.prifdmemaddr_17(\CPU|DP|prif.dmemaddr [17]),
	.prifdmemaddr_16(\CPU|DP|prif.dmemaddr [16]),
	.prifdmemaddr_19(\CPU|DP|prif.dmemaddr [19]),
	.prifdmemaddr_18(\CPU|DP|prif.dmemaddr [18]),
	.prifdmemaddr_25(\CPU|DP|prif.dmemaddr [25]),
	.prifdmemaddr_24(\CPU|DP|prif.dmemaddr [24]),
	.prifdmemaddr_27(\CPU|DP|prif.dmemaddr [27]),
	.prifdmemaddr_26(\CPU|DP|prif.dmemaddr [26]),
	.prifdmemstore_0(\CPU|DP|prif.dmemstore [0]),
	.prifdmemstore_1(\CPU|DP|prif.dmemstore [1]),
	.prifdmemstore_2(\CPU|DP|prif.dmemstore [2]),
	.prifdmemstore_3(\CPU|DP|prif.dmemstore [3]),
	.prifdmemstore_4(\CPU|DP|prif.dmemstore [4]),
	.prifdmemstore_5(\CPU|DP|prif.dmemstore [5]),
	.prifdmemstore_6(\CPU|DP|prif.dmemstore [6]),
	.prifdmemstore_7(\CPU|DP|prif.dmemstore [7]),
	.prifdmemstore_8(\CPU|DP|prif.dmemstore [8]),
	.prifdmemstore_9(\CPU|DP|prif.dmemstore [9]),
	.prifdmemstore_10(\CPU|DP|prif.dmemstore [10]),
	.prifdmemstore_11(\CPU|DP|prif.dmemstore [11]),
	.prifdmemstore_12(\CPU|DP|prif.dmemstore [12]),
	.prifdmemstore_13(\CPU|DP|prif.dmemstore [13]),
	.prifdmemstore_14(\CPU|DP|prif.dmemstore [14]),
	.prifdmemstore_15(\CPU|DP|prif.dmemstore [15]),
	.prifdmemstore_16(\CPU|DP|prif.dmemstore [16]),
	.prifdmemstore_17(\CPU|DP|prif.dmemstore [17]),
	.prifdmemstore_18(\CPU|DP|prif.dmemstore [18]),
	.prifdmemstore_19(\CPU|DP|prif.dmemstore [19]),
	.prifdmemstore_20(\CPU|DP|prif.dmemstore [20]),
	.prifdmemstore_21(\CPU|DP|prif.dmemstore [21]),
	.prifdmemstore_22(\CPU|DP|prif.dmemstore [22]),
	.prifdmemstore_23(\CPU|DP|prif.dmemstore [23]),
	.prifdmemstore_24(\CPU|DP|prif.dmemstore [24]),
	.prifdmemstore_25(\CPU|DP|prif.dmemstore [25]),
	.prifdmemstore_26(\CPU|DP|prif.dmemstore [26]),
	.prifdmemstore_27(\CPU|DP|prif.dmemstore [27]),
	.prifdmemstore_28(\CPU|DP|prif.dmemstore [28]),
	.prifdmemstore_29(\CPU|DP|prif.dmemstore [29]),
	.prifdmemstore_30(\CPU|DP|prif.dmemstore [30]),
	.prifdmemstore_31(\CPU|DP|prif.dmemstore [31]),
	.LessThan1(\RAM|LessThan1~0_combout ),
	.pc_3(\CPU|DP|pc [3]),
	.pc_2(\CPU|DP|pc [2]),
	.pc_5(\CPU|DP|pc [5]),
	.pc_4(\CPU|DP|pc [4]),
	.pc_7(\CPU|DP|pc [7]),
	.pc_6(\CPU|DP|pc [6]),
	.pc_9(\CPU|DP|pc [9]),
	.pc_8(\CPU|DP|pc [8]),
	.pc_11(\CPU|DP|pc [11]),
	.pc_10(\CPU|DP|pc [10]),
	.pc_13(\CPU|DP|pc [13]),
	.pc_12(\CPU|DP|pc [12]),
	.pc_15(\CPU|DP|pc [15]),
	.pc_14(\CPU|DP|pc [14]),
	.pc_23(\CPU|DP|pc [23]),
	.pc_22(\CPU|DP|pc [22]),
	.pc_21(\CPU|DP|pc [21]),
	.pc_29(\CPU|DP|pc [29]),
	.pc_28(\CPU|DP|pc [28]),
	.pc_31(\CPU|DP|pc [31]),
	.pc_30(\CPU|DP|pc [30]),
	.pc_20(\CPU|DP|pc [20]),
	.pc_17(\CPU|DP|pc [17]),
	.pc_16(\CPU|DP|pc [16]),
	.pc_19(\CPU|DP|pc [19]),
	.pc_18(\CPU|DP|pc [18]),
	.pc_25(\CPU|DP|pc [25]),
	.pc_24(\CPU|DP|pc [24]),
	.pc_27(\CPU|DP|pc [27]),
	.pc_26(\CPU|DP|pc [26]),
	.always0(\RAM|always0~21_combout ),
	.always1(\RAM|always1~0_combout ),
	.ramiframload_0(\RAM|ramif.ramload[0]~0_combout ),
	.ramiframload_1(\RAM|ramif.ramload[1]~1_combout ),
	.ramiframload_2(\RAM|ramif.ramload[2]~2_combout ),
	.ramiframload_3(\RAM|ramif.ramload[3]~3_combout ),
	.ramiframload_4(\RAM|ramif.ramload[4]~4_combout ),
	.ramiframload_5(\RAM|ramif.ramload[5]~5_combout ),
	.ramiframload_6(\RAM|ramif.ramload[6]~6_combout ),
	.ramiframload_7(\RAM|ramif.ramload[7]~7_combout ),
	.ramiframload_8(\RAM|ramif.ramload[8]~8_combout ),
	.ramiframload_9(\RAM|ramif.ramload[9]~9_combout ),
	.ramiframload_10(\RAM|ramif.ramload[10]~10_combout ),
	.ramiframload_11(\RAM|ramif.ramload[11]~11_combout ),
	.ramiframload_12(\RAM|ramif.ramload[12]~12_combout ),
	.ramiframload_13(\RAM|ramif.ramload[13]~13_combout ),
	.ramiframload_14(\RAM|ramif.ramload[14]~14_combout ),
	.ramiframload_15(\RAM|ramif.ramload[15]~15_combout ),
	.ramiframload_16(\RAM|ramif.ramload[16]~16_combout ),
	.ramiframload_17(\RAM|ramif.ramload[17]~17_combout ),
	.ramiframload_18(\RAM|ramif.ramload[18]~18_combout ),
	.ramiframload_19(\RAM|ramif.ramload[19]~19_combout ),
	.ramiframload_20(\RAM|ramif.ramload[20]~20_combout ),
	.ramiframload_21(\RAM|ramif.ramload[21]~21_combout ),
	.ramiframload_22(\RAM|ramif.ramload[22]~22_combout ),
	.ramiframload_23(\RAM|ramif.ramload[23]~23_combout ),
	.ramiframload_24(\RAM|ramif.ramload[24]~24_combout ),
	.ramiframload_25(\RAM|ramif.ramload[25]~25_combout ),
	.ramiframload_26(\RAM|ramif.ramload[26]~26_combout ),
	.ramiframload_27(\RAM|ramif.ramload[27]~27_combout ),
	.ramiframload_28(\RAM|ramif.ramload[28]~28_combout ),
	.ramiframload_29(\RAM|ramif.ramload[29]~29_combout ),
	.ramiframload_30(\RAM|ramif.ramload[30]~30_combout ),
	.ramiframload_31(\RAM|ramif.ramload[31]~31_combout ),
	.nRST(\nRST~input_o ),
	.CLK(\CPUCLK~clkctrl_outclk ),
	.nRST1(\nRST~inputclkctrl_outclk ),
	.dpifhalt(\CPU|DP|dpif.halt~q ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X60_Y29_N24
cycloneive_lcell_comb \ramaddr~0 (
// Equation(s):
// \ramaddr~0_combout  = (prifdmemwen & (((prifdmemaddr_1)))) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_1)) # (!prifdmemren & ((pc_1)))))

	.dataa(\CPU|DP|prif.dmemwen~q ),
	.datab(\CPU|DP|prif.dmemren~q ),
	.datac(\CPU|DP|prif.dmemaddr [1]),
	.datad(\CPU|DP|pc [1]),
	.cin(gnd),
	.combout(\ramaddr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~0 .lut_mask = 16'hF1E0;
defparam \ramaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N2
cycloneive_lcell_comb \ramaddr~1 (
// Equation(s):
// \ramaddr~1_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~0_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[1]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~0_combout ),
	.cin(gnd),
	.combout(\ramaddr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~1 .lut_mask = 16'hDD88;
defparam \ramaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N18
cycloneive_lcell_comb \ramaddr~2 (
// Equation(s):
// \ramaddr~2_combout  = (prifdmemwen & (((prifdmemaddr_0)))) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_0)) # (!prifdmemren & ((pc_0)))))

	.dataa(\CPU|DP|prif.dmemwen~q ),
	.datab(\CPU|DP|prif.dmemren~q ),
	.datac(\CPU|DP|prif.dmemaddr [0]),
	.datad(\CPU|DP|pc [0]),
	.cin(gnd),
	.combout(\ramaddr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~2 .lut_mask = 16'hF1E0;
defparam \ramaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N12
cycloneive_lcell_comb \ramaddr~3 (
// Equation(s):
// \ramaddr~3_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~2_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[0]~input_o ),
	.datad(\ramaddr~2_combout ),
	.cin(gnd),
	.combout(\ramaddr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~3 .lut_mask = 16'hF5A0;
defparam \ramaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N22
cycloneive_lcell_comb \ramaddr~4 (
// Equation(s):
// \ramaddr~4_combout  = (prifdmemwen & (((prifdmemaddr_3)))) # (!prifdmemwen & ((prifdmemren & ((prifdmemaddr_3))) # (!prifdmemren & (pc_3))))

	.dataa(\CPU|DP|prif.dmemwen~q ),
	.datab(\CPU|DP|pc [3]),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|prif.dmemaddr [3]),
	.cin(gnd),
	.combout(\ramaddr~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~4 .lut_mask = 16'hFE04;
defparam \ramaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N10
cycloneive_lcell_comb \ramaddr~5 (
// Equation(s):
// \ramaddr~5_combout  = (\syif.tbCTRL~input_o  & ((\syif.addr[3]~input_o ))) # (!\syif.tbCTRL~input_o  & (\ramaddr~4_combout ))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\ramaddr~4_combout ),
	.datad(\syif.addr[3]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~5 .lut_mask = 16'hFA50;
defparam \ramaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N6
cycloneive_lcell_comb \ramaddr~6 (
// Equation(s):
// \ramaddr~6_combout  = (prifdmemwen & (((prifdmemaddr_2)))) # (!prifdmemwen & ((prifdmemren & ((prifdmemaddr_2))) # (!prifdmemren & (pc_2))))

	.dataa(\CPU|DP|prif.dmemwen~q ),
	.datab(\CPU|DP|pc [2]),
	.datac(\CPU|DP|prif.dmemaddr [2]),
	.datad(\CPU|DP|prif.dmemren~q ),
	.cin(gnd),
	.combout(\ramaddr~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~6 .lut_mask = 16'hF0E4;
defparam \ramaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N16
cycloneive_lcell_comb \ramaddr~7 (
// Equation(s):
// \ramaddr~7_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[2]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~6_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(\syif.addr[2]~input_o ),
	.datac(gnd),
	.datad(\ramaddr~6_combout ),
	.cin(gnd),
	.combout(\ramaddr~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~7 .lut_mask = 16'hDD88;
defparam \ramaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N28
cycloneive_lcell_comb \ramaddr~8 (
// Equation(s):
// \ramaddr~8_combout  = (prifdmemwen & (prifdmemaddr_5)) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_5)) # (!prifdmemren & ((pc_5)))))

	.dataa(\CPU|DP|prif.dmemwen~q ),
	.datab(\CPU|DP|prif.dmemaddr [5]),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|pc [5]),
	.cin(gnd),
	.combout(\ramaddr~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~8 .lut_mask = 16'hCDC8;
defparam \ramaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N6
cycloneive_lcell_comb \ramaddr~9 (
// Equation(s):
// \ramaddr~9_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~8_combout )))

	.dataa(\syif.addr[5]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~8_combout ),
	.cin(gnd),
	.combout(\ramaddr~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~9 .lut_mask = 16'hAFA0;
defparam \ramaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N10
cycloneive_lcell_comb \ramaddr~10 (
// Equation(s):
// \ramaddr~10_combout  = (prifdmemwen & (((prifdmemaddr_4)))) # (!prifdmemwen & ((prifdmemren & ((prifdmemaddr_4))) # (!prifdmemren & (pc_4))))

	.dataa(\CPU|DP|prif.dmemwen~q ),
	.datab(\CPU|DP|pc [4]),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|prif.dmemaddr [4]),
	.cin(gnd),
	.combout(\ramaddr~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~10 .lut_mask = 16'hFE04;
defparam \ramaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N4
cycloneive_lcell_comb \ramaddr~11 (
// Equation(s):
// \ramaddr~11_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[4]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~10_combout )))

	.dataa(gnd),
	.datab(\syif.addr[4]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~10_combout ),
	.cin(gnd),
	.combout(\ramaddr~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~11 .lut_mask = 16'hCFC0;
defparam \ramaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N28
cycloneive_lcell_comb \ramaddr~12 (
// Equation(s):
// \ramaddr~12_combout  = (prifdmemwen & (prifdmemaddr_7)) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_7)) # (!prifdmemren & ((pc_7)))))

	.dataa(\CPU|DP|prif.dmemaddr [7]),
	.datab(\CPU|DP|pc [7]),
	.datac(\CPU|DP|prif.dmemwen~q ),
	.datad(\CPU|DP|prif.dmemren~q ),
	.cin(gnd),
	.combout(\ramaddr~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~12 .lut_mask = 16'hAAAC;
defparam \ramaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N22
cycloneive_lcell_comb \ramaddr~13 (
// Equation(s):
// \ramaddr~13_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~12_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[7]~input_o ),
	.datad(\ramaddr~12_combout ),
	.cin(gnd),
	.combout(\ramaddr~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~13 .lut_mask = 16'hF5A0;
defparam \ramaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N10
cycloneive_lcell_comb \ramaddr~14 (
// Equation(s):
// \ramaddr~14_combout  = (prifdmemwen & (((prifdmemaddr_6)))) # (!prifdmemwen & ((prifdmemren & ((prifdmemaddr_6))) # (!prifdmemren & (pc_6))))

	.dataa(\CPU|DP|pc [6]),
	.datab(\CPU|DP|prif.dmemaddr [6]),
	.datac(\CPU|DP|prif.dmemwen~q ),
	.datad(\CPU|DP|prif.dmemren~q ),
	.cin(gnd),
	.combout(\ramaddr~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~14 .lut_mask = 16'hCCCA;
defparam \ramaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N16
cycloneive_lcell_comb \ramaddr~15 (
// Equation(s):
// \ramaddr~15_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~14_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[6]~input_o ),
	.datad(\ramaddr~14_combout ),
	.cin(gnd),
	.combout(\ramaddr~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~15 .lut_mask = 16'hF5A0;
defparam \ramaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N24
cycloneive_lcell_comb \ramaddr~16 (
// Equation(s):
// \ramaddr~16_combout  = (prifdmemwen & (((prifdmemaddr_9)))) # (!prifdmemwen & ((prifdmemren & ((prifdmemaddr_9))) # (!prifdmemren & (pc_9))))

	.dataa(\CPU|DP|pc [9]),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|prif.dmemaddr [9]),
	.cin(gnd),
	.combout(\ramaddr~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~16 .lut_mask = 16'hFE02;
defparam \ramaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N26
cycloneive_lcell_comb \ramaddr~17 (
// Equation(s):
// \ramaddr~17_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~16_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[9]~input_o ),
	.datad(\ramaddr~16_combout ),
	.cin(gnd),
	.combout(\ramaddr~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~17 .lut_mask = 16'hF3C0;
defparam \ramaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N18
cycloneive_lcell_comb \ramaddr~18 (
// Equation(s):
// \ramaddr~18_combout  = (prifdmemwen & (prifdmemaddr_8)) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_8)) # (!prifdmemren & ((pc_8)))))

	.dataa(\CPU|DP|prif.dmemaddr [8]),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|pc [8]),
	.cin(gnd),
	.combout(\ramaddr~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~18 .lut_mask = 16'hABA8;
defparam \ramaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N0
cycloneive_lcell_comb \ramaddr~19 (
// Equation(s):
// \ramaddr~19_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~18_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[8]~input_o ),
	.datad(\ramaddr~18_combout ),
	.cin(gnd),
	.combout(\ramaddr~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~19 .lut_mask = 16'hF3C0;
defparam \ramaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N10
cycloneive_lcell_comb \ramaddr~20 (
// Equation(s):
// \ramaddr~20_combout  = (prifdmemren & (prifdmemaddr_11)) # (!prifdmemren & ((prifdmemwen & (prifdmemaddr_11)) # (!prifdmemwen & ((pc_11)))))

	.dataa(\CPU|DP|prif.dmemaddr [11]),
	.datab(\CPU|DP|prif.dmemren~q ),
	.datac(\CPU|DP|pc [11]),
	.datad(\CPU|DP|prif.dmemwen~q ),
	.cin(gnd),
	.combout(\ramaddr~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~20 .lut_mask = 16'hAAB8;
defparam \ramaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N28
cycloneive_lcell_comb \ramaddr~21 (
// Equation(s):
// \ramaddr~21_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~20_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[11]~input_o ),
	.datad(\ramaddr~20_combout ),
	.cin(gnd),
	.combout(\ramaddr~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~21 .lut_mask = 16'hF3C0;
defparam \ramaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N20
cycloneive_lcell_comb \ramaddr~22 (
// Equation(s):
// \ramaddr~22_combout  = (prifdmemren & (prifdmemaddr_10)) # (!prifdmemren & ((prifdmemwen & (prifdmemaddr_10)) # (!prifdmemwen & ((pc_10)))))

	.dataa(\CPU|DP|prif.dmemaddr [10]),
	.datab(\CPU|DP|prif.dmemren~q ),
	.datac(\CPU|DP|pc [10]),
	.datad(\CPU|DP|prif.dmemwen~q ),
	.cin(gnd),
	.combout(\ramaddr~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~22 .lut_mask = 16'hAAB8;
defparam \ramaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N2
cycloneive_lcell_comb \ramaddr~23 (
// Equation(s):
// \ramaddr~23_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~22_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[10]~input_o ),
	.datad(\ramaddr~22_combout ),
	.cin(gnd),
	.combout(\ramaddr~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~23 .lut_mask = 16'hF3C0;
defparam \ramaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N2
cycloneive_lcell_comb \ramaddr~24 (
// Equation(s):
// \ramaddr~24_combout  = (prifdmemwen & (prifdmemaddr_13)) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_13)) # (!prifdmemren & ((pc_13)))))

	.dataa(\CPU|DP|prif.dmemaddr [13]),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|pc [13]),
	.cin(gnd),
	.combout(\ramaddr~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~24 .lut_mask = 16'hABA8;
defparam \ramaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N4
cycloneive_lcell_comb \ramaddr~25 (
// Equation(s):
// \ramaddr~25_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[13]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~24_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[13]~input_o ),
	.datad(\ramaddr~24_combout ),
	.cin(gnd),
	.combout(\ramaddr~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~25 .lut_mask = 16'hF3C0;
defparam \ramaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N28
cycloneive_lcell_comb \ramaddr~26 (
// Equation(s):
// \ramaddr~26_combout  = (prifdmemwen & (prifdmemaddr_12)) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_12)) # (!prifdmemren & ((pc_12)))))

	.dataa(\CPU|DP|prif.dmemaddr [12]),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|pc [12]),
	.cin(gnd),
	.combout(\ramaddr~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~26 .lut_mask = 16'hABA8;
defparam \ramaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N6
cycloneive_lcell_comb \ramaddr~27 (
// Equation(s):
// \ramaddr~27_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~26_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[12]~input_o ),
	.datad(\ramaddr~26_combout ),
	.cin(gnd),
	.combout(\ramaddr~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~27 .lut_mask = 16'hF3C0;
defparam \ramaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N24
cycloneive_lcell_comb \ramaddr~28 (
// Equation(s):
// \ramaddr~28_combout  = (prifdmemwen & (((prifdmemaddr_15)))) # (!prifdmemwen & ((prifdmemren & ((prifdmemaddr_15))) # (!prifdmemren & (pc_15))))

	.dataa(\CPU|DP|pc [15]),
	.datab(\CPU|DP|prif.dmemaddr [15]),
	.datac(\CPU|DP|prif.dmemwen~q ),
	.datad(\CPU|DP|prif.dmemren~q ),
	.cin(gnd),
	.combout(\ramaddr~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~28 .lut_mask = 16'hCCCA;
defparam \ramaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N26
cycloneive_lcell_comb \ramaddr~29 (
// Equation(s):
// \ramaddr~29_combout  = (\syif.tbCTRL~input_o  & (!\syif.addr[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((!\ramaddr~28_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[15]~input_o ),
	.datad(\ramaddr~28_combout ),
	.cin(gnd),
	.combout(\ramaddr~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29 .lut_mask = 16'h0C3F;
defparam \ramaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N16
cycloneive_lcell_comb \ramaddr~30 (
// Equation(s):
// \ramaddr~30_combout  = (prifdmemwen & (prifdmemaddr_14)) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_14)) # (!prifdmemren & ((pc_14)))))

	.dataa(\CPU|DP|prif.dmemaddr [14]),
	.datab(\CPU|DP|pc [14]),
	.datac(\CPU|DP|prif.dmemwen~q ),
	.datad(\CPU|DP|prif.dmemren~q ),
	.cin(gnd),
	.combout(\ramaddr~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~30 .lut_mask = 16'hAAAC;
defparam \ramaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N2
cycloneive_lcell_comb \ramaddr~31 (
// Equation(s):
// \ramaddr~31_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~30_combout )))

	.dataa(gnd),
	.datab(\syif.addr[14]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~30_combout ),
	.cin(gnd),
	.combout(\ramaddr~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~31 .lut_mask = 16'hCFC0;
defparam \ramaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N28
cycloneive_lcell_comb \ramaddr~32 (
// Equation(s):
// \ramaddr~32_combout  = (prifdmemren & (((prifdmemaddr_23)))) # (!prifdmemren & ((prifdmemwen & ((prifdmemaddr_23))) # (!prifdmemwen & (pc_23))))

	.dataa(\CPU|DP|prif.dmemren~q ),
	.datab(\CPU|DP|pc [23]),
	.datac(\CPU|DP|prif.dmemaddr [23]),
	.datad(\CPU|DP|prif.dmemwen~q ),
	.cin(gnd),
	.combout(\ramaddr~32_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~32 .lut_mask = 16'hF0E4;
defparam \ramaddr~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N6
cycloneive_lcell_comb \ramaddr~33 (
// Equation(s):
// \ramaddr~33_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~32_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[23]~input_o ),
	.datad(\ramaddr~32_combout ),
	.cin(gnd),
	.combout(\ramaddr~33_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~33 .lut_mask = 16'hF3C0;
defparam \ramaddr~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N18
cycloneive_lcell_comb \ramaddr~34 (
// Equation(s):
// \ramaddr~34_combout  = (prifdmemwen & (prifdmemaddr_22)) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_22)) # (!prifdmemren & ((pc_22)))))

	.dataa(\CPU|DP|prif.dmemwen~q ),
	.datab(\CPU|DP|prif.dmemaddr [22]),
	.datac(\CPU|DP|pc [22]),
	.datad(\CPU|DP|prif.dmemren~q ),
	.cin(gnd),
	.combout(\ramaddr~34_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~34 .lut_mask = 16'hCCD8;
defparam \ramaddr~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N12
cycloneive_lcell_comb \ramaddr~35 (
// Equation(s):
// \ramaddr~35_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[22]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~34_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[22]~input_o ),
	.datad(\ramaddr~34_combout ),
	.cin(gnd),
	.combout(\ramaddr~35_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~35 .lut_mask = 16'hF3C0;
defparam \ramaddr~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N22
cycloneive_lcell_comb \ramWEN~0 (
// Equation(s):
// \ramWEN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.WEN~input_o )) # (!\syif.tbCTRL~input_o  & ((!prifdmemwen)))

	.dataa(\syif.WEN~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|prif.dmemwen~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramWEN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramWEN~0 .lut_mask = 16'h4747;
defparam \ramWEN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N4
cycloneive_lcell_comb \ramREN~0 (
// Equation(s):
// \ramREN~0_combout  = (\syif.tbCTRL~input_o  & (!\syif.REN~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemwen)))

	.dataa(\syif.REN~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|prif.dmemwen~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramREN~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramREN~0 .lut_mask = 16'h7474;
defparam \ramREN~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N28
cycloneive_lcell_comb \ramaddr~36 (
// Equation(s):
// \ramaddr~36_combout  = (prifdmemwen & (((prifdmemaddr_21)))) # (!prifdmemwen & ((prifdmemren & ((prifdmemaddr_21))) # (!prifdmemren & (pc_21))))

	.dataa(\CPU|DP|pc [21]),
	.datab(\CPU|DP|prif.dmemaddr [21]),
	.datac(\CPU|DP|prif.dmemwen~q ),
	.datad(\CPU|DP|prif.dmemren~q ),
	.cin(gnd),
	.combout(\ramaddr~36_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~36 .lut_mask = 16'hCCCA;
defparam \ramaddr~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N10
cycloneive_lcell_comb \ramaddr~37 (
// Equation(s):
// \ramaddr~37_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[21]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~36_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[21]~input_o ),
	.datad(\ramaddr~36_combout ),
	.cin(gnd),
	.combout(\ramaddr~37_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~37 .lut_mask = 16'hF3C0;
defparam \ramaddr~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N12
cycloneive_lcell_comb \ramaddr~38 (
// Equation(s):
// \ramaddr~38_combout  = (prifdmemren & (((prifdmemaddr_29)))) # (!prifdmemren & ((prifdmemwen & ((prifdmemaddr_29))) # (!prifdmemwen & (pc_29))))

	.dataa(\CPU|DP|prif.dmemren~q ),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|pc [29]),
	.datad(\CPU|DP|prif.dmemaddr [29]),
	.cin(gnd),
	.combout(\ramaddr~38_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~38 .lut_mask = 16'hFE10;
defparam \ramaddr~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N6
cycloneive_lcell_comb \ramaddr~39 (
// Equation(s):
// \ramaddr~39_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[29]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~38_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[29]~input_o ),
	.datad(\ramaddr~38_combout ),
	.cin(gnd),
	.combout(\ramaddr~39_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~39 .lut_mask = 16'hF3C0;
defparam \ramaddr~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N10
cycloneive_lcell_comb \ramaddr~40 (
// Equation(s):
// \ramaddr~40_combout  = (prifdmemren & (((prifdmemaddr_28)))) # (!prifdmemren & ((prifdmemwen & ((prifdmemaddr_28))) # (!prifdmemwen & (pc_28))))

	.dataa(\CPU|DP|prif.dmemren~q ),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|pc [28]),
	.datad(\CPU|DP|prif.dmemaddr [28]),
	.cin(gnd),
	.combout(\ramaddr~40_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~40 .lut_mask = 16'hFE10;
defparam \ramaddr~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N4
cycloneive_lcell_comb \ramaddr~41 (
// Equation(s):
// \ramaddr~41_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~40_combout )))

	.dataa(\syif.addr[28]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~40_combout ),
	.cin(gnd),
	.combout(\ramaddr~41_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~41 .lut_mask = 16'hBB88;
defparam \ramaddr~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N18
cycloneive_lcell_comb \ramaddr~42 (
// Equation(s):
// \ramaddr~42_combout  = (prifdmemren & (((prifdmemaddr_31)))) # (!prifdmemren & ((prifdmemwen & (prifdmemaddr_31)) # (!prifdmemwen & ((pc_31)))))

	.dataa(\CPU|DP|prif.dmemren~q ),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|prif.dmemaddr [31]),
	.datad(\CPU|DP|pc [31]),
	.cin(gnd),
	.combout(\ramaddr~42_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~42 .lut_mask = 16'hF1E0;
defparam \ramaddr~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N0
cycloneive_lcell_comb \ramaddr~43 (
// Equation(s):
// \ramaddr~43_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~42_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[31]~input_o ),
	.datad(\ramaddr~42_combout ),
	.cin(gnd),
	.combout(\ramaddr~43_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~43 .lut_mask = 16'hF3C0;
defparam \ramaddr~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N20
cycloneive_lcell_comb \ramaddr~44 (
// Equation(s):
// \ramaddr~44_combout  = (prifdmemren & (((prifdmemaddr_30)))) # (!prifdmemren & ((prifdmemwen & (prifdmemaddr_30)) # (!prifdmemwen & ((pc_30)))))

	.dataa(\CPU|DP|prif.dmemren~q ),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|prif.dmemaddr [30]),
	.datad(\CPU|DP|pc [30]),
	.cin(gnd),
	.combout(\ramaddr~44_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~44 .lut_mask = 16'hF1E0;
defparam \ramaddr~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N22
cycloneive_lcell_comb \ramaddr~45 (
// Equation(s):
// \ramaddr~45_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[30]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~44_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[30]~input_o ),
	.datad(\ramaddr~44_combout ),
	.cin(gnd),
	.combout(\ramaddr~45_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~45 .lut_mask = 16'hF3C0;
defparam \ramaddr~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N16
cycloneive_lcell_comb \ramaddr~46 (
// Equation(s):
// \ramaddr~46_combout  = (prifdmemwen & (prifdmemaddr_20)) # (!prifdmemwen & ((prifdmemren & (prifdmemaddr_20)) # (!prifdmemren & ((pc_20)))))

	.dataa(\CPU|DP|prif.dmemwen~q ),
	.datab(\CPU|DP|prif.dmemaddr [20]),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|pc [20]),
	.cin(gnd),
	.combout(\ramaddr~46_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~46 .lut_mask = 16'hCDC8;
defparam \ramaddr~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N22
cycloneive_lcell_comb \ramaddr~47 (
// Equation(s):
// \ramaddr~47_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~46_combout )))

	.dataa(gnd),
	.datab(\syif.addr[20]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~46_combout ),
	.cin(gnd),
	.combout(\ramaddr~47_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~47 .lut_mask = 16'hCFC0;
defparam \ramaddr~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N6
cycloneive_lcell_comb \ramaddr~48 (
// Equation(s):
// \ramaddr~48_combout  = (prifdmemren & (prifdmemaddr_17)) # (!prifdmemren & ((prifdmemwen & (prifdmemaddr_17)) # (!prifdmemwen & ((pc_17)))))

	.dataa(\CPU|DP|prif.dmemren~q ),
	.datab(\CPU|DP|prif.dmemaddr [17]),
	.datac(\CPU|DP|pc [17]),
	.datad(\CPU|DP|prif.dmemwen~q ),
	.cin(gnd),
	.combout(\ramaddr~48_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~48 .lut_mask = 16'hCCD8;
defparam \ramaddr~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N16
cycloneive_lcell_comb \ramaddr~49 (
// Equation(s):
// \ramaddr~49_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[17]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~48_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[17]~input_o ),
	.datad(\ramaddr~48_combout ),
	.cin(gnd),
	.combout(\ramaddr~49_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~49 .lut_mask = 16'hF3C0;
defparam \ramaddr~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N24
cycloneive_lcell_comb \ramaddr~50 (
// Equation(s):
// \ramaddr~50_combout  = (prifdmemren & (prifdmemaddr_16)) # (!prifdmemren & ((prifdmemwen & (prifdmemaddr_16)) # (!prifdmemwen & ((pc_16)))))

	.dataa(\CPU|DP|prif.dmemaddr [16]),
	.datab(\CPU|DP|pc [16]),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|prif.dmemwen~q ),
	.cin(gnd),
	.combout(\ramaddr~50_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~50 .lut_mask = 16'hAAAC;
defparam \ramaddr~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N30
cycloneive_lcell_comb \ramaddr~51 (
// Equation(s):
// \ramaddr~51_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[16]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~50_combout )))

	.dataa(\syif.addr[16]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\ramaddr~50_combout ),
	.cin(gnd),
	.combout(\ramaddr~51_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~51 .lut_mask = 16'hBB88;
defparam \ramaddr~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N10
cycloneive_lcell_comb \ramaddr~52 (
// Equation(s):
// \ramaddr~52_combout  = (prifdmemren & (((prifdmemaddr_19)))) # (!prifdmemren & ((prifdmemwen & ((prifdmemaddr_19))) # (!prifdmemwen & (pc_19))))

	.dataa(\CPU|DP|pc [19]),
	.datab(\CPU|DP|prif.dmemaddr [19]),
	.datac(\CPU|DP|prif.dmemren~q ),
	.datad(\CPU|DP|prif.dmemwen~q ),
	.cin(gnd),
	.combout(\ramaddr~52_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~52 .lut_mask = 16'hCCCA;
defparam \ramaddr~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N28
cycloneive_lcell_comb \ramaddr~53 (
// Equation(s):
// \ramaddr~53_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~52_combout )))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.addr[19]~input_o ),
	.datad(\ramaddr~52_combout ),
	.cin(gnd),
	.combout(\ramaddr~53_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~53 .lut_mask = 16'hF3C0;
defparam \ramaddr~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N20
cycloneive_lcell_comb \ramaddr~54 (
// Equation(s):
// \ramaddr~54_combout  = (prifdmemren & (((prifdmemaddr_18)))) # (!prifdmemren & ((prifdmemwen & ((prifdmemaddr_18))) # (!prifdmemwen & (pc_18))))

	.dataa(\CPU|DP|pc [18]),
	.datab(\CPU|DP|prif.dmemren~q ),
	.datac(\CPU|DP|prif.dmemwen~q ),
	.datad(\CPU|DP|prif.dmemaddr [18]),
	.cin(gnd),
	.combout(\ramaddr~54_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~54 .lut_mask = 16'hFE02;
defparam \ramaddr~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N22
cycloneive_lcell_comb \ramaddr~55 (
// Equation(s):
// \ramaddr~55_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~54_combout )))

	.dataa(gnd),
	.datab(\syif.addr[18]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~54_combout ),
	.cin(gnd),
	.combout(\ramaddr~55_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~55 .lut_mask = 16'hCFC0;
defparam \ramaddr~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N30
cycloneive_lcell_comb \ramaddr~56 (
// Equation(s):
// \ramaddr~56_combout  = (prifdmemren & (prifdmemaddr_25)) # (!prifdmemren & ((prifdmemwen & (prifdmemaddr_25)) # (!prifdmemwen & ((pc_25)))))

	.dataa(\CPU|DP|prif.dmemaddr [25]),
	.datab(\CPU|DP|prif.dmemren~q ),
	.datac(\CPU|DP|prif.dmemwen~q ),
	.datad(\CPU|DP|pc [25]),
	.cin(gnd),
	.combout(\ramaddr~56_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~56 .lut_mask = 16'hABA8;
defparam \ramaddr~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N16
cycloneive_lcell_comb \ramaddr~57 (
// Equation(s):
// \ramaddr~57_combout  = (\syif.tbCTRL~input_o  & ((\syif.addr[25]~input_o ))) # (!\syif.tbCTRL~input_o  & (\ramaddr~56_combout ))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\ramaddr~56_combout ),
	.datad(\syif.addr[25]~input_o ),
	.cin(gnd),
	.combout(\ramaddr~57_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~57 .lut_mask = 16'hFC30;
defparam \ramaddr~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N28
cycloneive_lcell_comb \ramaddr~58 (
// Equation(s):
// \ramaddr~58_combout  = (prifdmemwen & (((prifdmemaddr_24)))) # (!prifdmemwen & ((prifdmemren & ((prifdmemaddr_24))) # (!prifdmemren & (pc_24))))

	.dataa(\CPU|DP|pc [24]),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|prif.dmemaddr [24]),
	.datad(\CPU|DP|prif.dmemren~q ),
	.cin(gnd),
	.combout(\ramaddr~58_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~58 .lut_mask = 16'hF0E2;
defparam \ramaddr~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N26
cycloneive_lcell_comb \ramaddr~59 (
// Equation(s):
// \ramaddr~59_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~58_combout )))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\syif.addr[24]~input_o ),
	.datad(\ramaddr~58_combout ),
	.cin(gnd),
	.combout(\ramaddr~59_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~59 .lut_mask = 16'hF5A0;
defparam \ramaddr~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N24
cycloneive_lcell_comb \ramaddr~60 (
// Equation(s):
// \ramaddr~60_combout  = (prifdmemren & (((prifdmemaddr_27)))) # (!prifdmemren & ((prifdmemwen & ((prifdmemaddr_27))) # (!prifdmemwen & (pc_27))))

	.dataa(\CPU|DP|prif.dmemren~q ),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|pc [27]),
	.datad(\CPU|DP|prif.dmemaddr [27]),
	.cin(gnd),
	.combout(\ramaddr~60_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~60 .lut_mask = 16'hFE10;
defparam \ramaddr~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N20
cycloneive_lcell_comb \ramaddr~61 (
// Equation(s):
// \ramaddr~61_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~60_combout )))

	.dataa(gnd),
	.datab(\syif.addr[27]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~60_combout ),
	.cin(gnd),
	.combout(\ramaddr~61_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~61 .lut_mask = 16'hCFC0;
defparam \ramaddr~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N2
cycloneive_lcell_comb \ramaddr~62 (
// Equation(s):
// \ramaddr~62_combout  = (prifdmemren & (((prifdmemaddr_26)))) # (!prifdmemren & ((prifdmemwen & (prifdmemaddr_26)) # (!prifdmemwen & ((pc_26)))))

	.dataa(\CPU|DP|prif.dmemren~q ),
	.datab(\CPU|DP|prif.dmemwen~q ),
	.datac(\CPU|DP|prif.dmemaddr [26]),
	.datad(\CPU|DP|pc [26]),
	.cin(gnd),
	.combout(\ramaddr~62_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~62 .lut_mask = 16'hF1E0;
defparam \ramaddr~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N6
cycloneive_lcell_comb \ramaddr~63 (
// Equation(s):
// \ramaddr~63_combout  = (\syif.tbCTRL~input_o  & (\syif.addr[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((\ramaddr~62_combout )))

	.dataa(gnd),
	.datab(\syif.addr[26]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\ramaddr~62_combout ),
	.cin(gnd),
	.combout(\ramaddr~63_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~63 .lut_mask = 16'hCFC0;
defparam \ramaddr~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y72_N7
dffeas CPUCLK(
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\CPUCLK~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\CPUCLK~q ),
	.prn(vcc));
// synopsys translate_off
defparam CPUCLK.is_wysiwyg = "true";
defparam CPUCLK.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N12
cycloneive_lcell_comb \ramstore~0 (
// Equation(s):
// \ramstore~0_combout  = (\syif.tbCTRL~input_o  & (\syif.store[0]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_0)))

	.dataa(\syif.store[0]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [0]),
	.cin(gnd),
	.combout(\ramstore~0_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~0 .lut_mask = 16'hAFA0;
defparam \ramstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N14
cycloneive_lcell_comb \ramstore~1 (
// Equation(s):
// \ramstore~1_combout  = (\syif.tbCTRL~input_o  & (\syif.store[1]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_1)))

	.dataa(\syif.store[1]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [1]),
	.cin(gnd),
	.combout(\ramstore~1_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~1 .lut_mask = 16'hAFA0;
defparam \ramstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y23_N30
cycloneive_lcell_comb \ramstore~2 (
// Equation(s):
// \ramstore~2_combout  = (\syif.tbCTRL~input_o  & (\syif.store[2]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_2)))

	.dataa(\syif.store[2]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [2]),
	.cin(gnd),
	.combout(\ramstore~2_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~2 .lut_mask = 16'hAFA0;
defparam \ramstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y22_N28
cycloneive_lcell_comb \ramstore~3 (
// Equation(s):
// \ramstore~3_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[3]~input_o ))) # (!\syif.tbCTRL~input_o  & (prifdmemstore_3))

	.dataa(\syif.tbCTRL~input_o ),
	.datab(gnd),
	.datac(\CPU|DP|prif.dmemstore [3]),
	.datad(\syif.store[3]~input_o ),
	.cin(gnd),
	.combout(\ramstore~3_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~3 .lut_mask = 16'hFA50;
defparam \ramstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N0
cycloneive_lcell_comb \ramstore~4 (
// Equation(s):
// \ramstore~4_combout  = (\syif.tbCTRL~input_o  & (\syif.store[4]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_4)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[4]~input_o ),
	.datad(\CPU|DP|prif.dmemstore [4]),
	.cin(gnd),
	.combout(\ramstore~4_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~4 .lut_mask = 16'hF3C0;
defparam \ramstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N22
cycloneive_lcell_comb \ramstore~5 (
// Equation(s):
// \ramstore~5_combout  = (\syif.tbCTRL~input_o  & (\syif.store[5]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_5)))

	.dataa(\syif.store[5]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [5]),
	.cin(gnd),
	.combout(\ramstore~5_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~5 .lut_mask = 16'hAFA0;
defparam \ramstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N8
cycloneive_lcell_comb \ramstore~6 (
// Equation(s):
// \ramstore~6_combout  = (\syif.tbCTRL~input_o  & (\syif.store[6]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_6)))

	.dataa(gnd),
	.datab(\syif.store[6]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [6]),
	.cin(gnd),
	.combout(\ramstore~6_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~6 .lut_mask = 16'hCFC0;
defparam \ramstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N26
cycloneive_lcell_comb \ramstore~7 (
// Equation(s):
// \ramstore~7_combout  = (\syif.tbCTRL~input_o  & (\syif.store[7]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_7)))

	.dataa(gnd),
	.datab(\syif.store[7]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [7]),
	.cin(gnd),
	.combout(\ramstore~7_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~7 .lut_mask = 16'hCFC0;
defparam \ramstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N30
cycloneive_lcell_comb \ramstore~8 (
// Equation(s):
// \ramstore~8_combout  = (\syif.tbCTRL~input_o  & (\syif.store[8]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_8)))

	.dataa(gnd),
	.datab(\syif.store[8]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [8]),
	.cin(gnd),
	.combout(\ramstore~8_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~8 .lut_mask = 16'hCFC0;
defparam \ramstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N0
cycloneive_lcell_comb \ramstore~9 (
// Equation(s):
// \ramstore~9_combout  = (\syif.tbCTRL~input_o  & (\syif.store[9]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_9)))

	.dataa(\syif.store[9]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [9]),
	.cin(gnd),
	.combout(\ramstore~9_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~9 .lut_mask = 16'hAFA0;
defparam \ramstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N8
cycloneive_lcell_comb \ramstore~10 (
// Equation(s):
// \ramstore~10_combout  = (\syif.tbCTRL~input_o  & (\syif.store[10]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_10)))

	.dataa(\syif.store[10]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [10]),
	.cin(gnd),
	.combout(\ramstore~10_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~10 .lut_mask = 16'hAFA0;
defparam \ramstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N22
cycloneive_lcell_comb \ramstore~11 (
// Equation(s):
// \ramstore~11_combout  = (\syif.tbCTRL~input_o  & (\syif.store[11]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_11)))

	.dataa(gnd),
	.datab(\syif.store[11]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [11]),
	.cin(gnd),
	.combout(\ramstore~11_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~11 .lut_mask = 16'hCFC0;
defparam \ramstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N4
cycloneive_lcell_comb \ramstore~12 (
// Equation(s):
// \ramstore~12_combout  = (\syif.tbCTRL~input_o  & (\syif.store[12]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_12)))

	.dataa(gnd),
	.datab(\syif.store[12]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [12]),
	.cin(gnd),
	.combout(\ramstore~12_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~12 .lut_mask = 16'hCFC0;
defparam \ramstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N28
cycloneive_lcell_comb \ramstore~13 (
// Equation(s):
// \ramstore~13_combout  = (\syif.tbCTRL~input_o  & (\syif.store[13]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_13)))

	.dataa(gnd),
	.datab(\syif.store[13]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [13]),
	.cin(gnd),
	.combout(\ramstore~13_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~13 .lut_mask = 16'hCFC0;
defparam \ramstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N30
cycloneive_lcell_comb \ramstore~14 (
// Equation(s):
// \ramstore~14_combout  = (\syif.tbCTRL~input_o  & (\syif.store[14]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_14)))

	.dataa(gnd),
	.datab(\syif.store[14]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [14]),
	.cin(gnd),
	.combout(\ramstore~14_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~14 .lut_mask = 16'hCFC0;
defparam \ramstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N0
cycloneive_lcell_comb \ramstore~15 (
// Equation(s):
// \ramstore~15_combout  = (\syif.tbCTRL~input_o  & (\syif.store[15]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_15)))

	.dataa(\syif.store[15]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [15]),
	.cin(gnd),
	.combout(\ramstore~15_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~15 .lut_mask = 16'hAFA0;
defparam \ramstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N14
cycloneive_lcell_comb \ramstore~16 (
// Equation(s):
// \ramstore~16_combout  = (\syif.tbCTRL~input_o  & (\syif.store[16]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_16)))

	.dataa(gnd),
	.datab(\syif.store[16]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [16]),
	.cin(gnd),
	.combout(\ramstore~16_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~16 .lut_mask = 16'hCFC0;
defparam \ramstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N16
cycloneive_lcell_comb \ramstore~17 (
// Equation(s):
// \ramstore~17_combout  = (\syif.tbCTRL~input_o  & (\syif.store[17]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_17)))

	.dataa(gnd),
	.datab(\syif.store[17]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [17]),
	.cin(gnd),
	.combout(\ramstore~17_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~17 .lut_mask = 16'hCFC0;
defparam \ramstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N26
cycloneive_lcell_comb \ramstore~18 (
// Equation(s):
// \ramstore~18_combout  = (\syif.tbCTRL~input_o  & (\syif.store[18]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_18)))

	.dataa(\syif.store[18]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [18]),
	.cin(gnd),
	.combout(\ramstore~18_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~18 .lut_mask = 16'hAFA0;
defparam \ramstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N14
cycloneive_lcell_comb \ramstore~19 (
// Equation(s):
// \ramstore~19_combout  = (\syif.tbCTRL~input_o  & (\syif.store[19]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_19)))

	.dataa(\syif.store[19]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [19]),
	.cin(gnd),
	.combout(\ramstore~19_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~19 .lut_mask = 16'hAFA0;
defparam \ramstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N24
cycloneive_lcell_comb \ramstore~20 (
// Equation(s):
// \ramstore~20_combout  = (\syif.tbCTRL~input_o  & (\syif.store[20]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_20)))

	.dataa(gnd),
	.datab(\syif.store[20]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [20]),
	.cin(gnd),
	.combout(\ramstore~20_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~20 .lut_mask = 16'hCFC0;
defparam \ramstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N30
cycloneive_lcell_comb \ramstore~21 (
// Equation(s):
// \ramstore~21_combout  = (\syif.tbCTRL~input_o  & (\syif.store[21]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_21)))

	.dataa(gnd),
	.datab(\syif.store[21]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [21]),
	.cin(gnd),
	.combout(\ramstore~21_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~21 .lut_mask = 16'hCFC0;
defparam \ramstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N22
cycloneive_lcell_comb \ramstore~22 (
// Equation(s):
// \ramstore~22_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[22]~input_o ))) # (!\syif.tbCTRL~input_o  & (prifdmemstore_22))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\CPU|DP|prif.dmemstore [22]),
	.datad(\syif.store[22]~input_o ),
	.cin(gnd),
	.combout(\ramstore~22_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~22 .lut_mask = 16'hFC30;
defparam \ramstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N8
cycloneive_lcell_comb \ramstore~23 (
// Equation(s):
// \ramstore~23_combout  = (\syif.tbCTRL~input_o  & (\syif.store[23]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_23)))

	.dataa(\syif.store[23]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [23]),
	.cin(gnd),
	.combout(\ramstore~23_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~23 .lut_mask = 16'hAFA0;
defparam \ramstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N8
cycloneive_lcell_comb \ramstore~24 (
// Equation(s):
// \ramstore~24_combout  = (\syif.tbCTRL~input_o  & (\syif.store[24]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_24)))

	.dataa(\syif.store[24]~input_o ),
	.datab(\syif.tbCTRL~input_o ),
	.datac(gnd),
	.datad(\CPU|DP|prif.dmemstore [24]),
	.cin(gnd),
	.combout(\ramstore~24_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~24 .lut_mask = 16'hBB88;
defparam \ramstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N18
cycloneive_lcell_comb \ramstore~25 (
// Equation(s):
// \ramstore~25_combout  = (\syif.tbCTRL~input_o  & (\syif.store[25]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_25)))

	.dataa(\syif.store[25]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [25]),
	.cin(gnd),
	.combout(\ramstore~25_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~25 .lut_mask = 16'hAFA0;
defparam \ramstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N28
cycloneive_lcell_comb \ramstore~26 (
// Equation(s):
// \ramstore~26_combout  = (\syif.tbCTRL~input_o  & (\syif.store[26]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_26)))

	.dataa(gnd),
	.datab(\syif.store[26]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [26]),
	.cin(gnd),
	.combout(\ramstore~26_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~26 .lut_mask = 16'hCFC0;
defparam \ramstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N28
cycloneive_lcell_comb \ramstore~27 (
// Equation(s):
// \ramstore~27_combout  = (\syif.tbCTRL~input_o  & (\syif.store[27]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_27)))

	.dataa(gnd),
	.datab(\syif.tbCTRL~input_o ),
	.datac(\syif.store[27]~input_o ),
	.datad(\CPU|DP|prif.dmemstore [27]),
	.cin(gnd),
	.combout(\ramstore~27_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~27 .lut_mask = 16'hF3C0;
defparam \ramstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N14
cycloneive_lcell_comb \ramstore~28 (
// Equation(s):
// \ramstore~28_combout  = (\syif.tbCTRL~input_o  & (\syif.store[28]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_28)))

	.dataa(gnd),
	.datab(\syif.store[28]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [28]),
	.cin(gnd),
	.combout(\ramstore~28_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~28 .lut_mask = 16'hCFC0;
defparam \ramstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N22
cycloneive_lcell_comb \ramstore~29 (
// Equation(s):
// \ramstore~29_combout  = (\syif.tbCTRL~input_o  & (\syif.store[29]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_29)))

	.dataa(\syif.store[29]~input_o ),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [29]),
	.cin(gnd),
	.combout(\ramstore~29_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~29 .lut_mask = 16'hAFA0;
defparam \ramstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N2
cycloneive_lcell_comb \ramstore~30 (
// Equation(s):
// \ramstore~30_combout  = (\syif.tbCTRL~input_o  & ((\syif.store[30]~input_o ))) # (!\syif.tbCTRL~input_o  & (prifdmemstore_30))

	.dataa(\CPU|DP|prif.dmemstore [30]),
	.datab(gnd),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\syif.store[30]~input_o ),
	.cin(gnd),
	.combout(\ramstore~30_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~30 .lut_mask = 16'hFA0A;
defparam \ramstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y21_N0
cycloneive_lcell_comb \ramstore~31 (
// Equation(s):
// \ramstore~31_combout  = (\syif.tbCTRL~input_o  & (\syif.store[31]~input_o )) # (!\syif.tbCTRL~input_o  & ((prifdmemstore_31)))

	.dataa(gnd),
	.datab(\syif.store[31]~input_o ),
	.datac(\syif.tbCTRL~input_o ),
	.datad(\CPU|DP|prif.dmemstore [31]),
	.cin(gnd),
	.combout(\ramstore~31_combout ),
	.cout());
// synopsys translate_off
defparam \ramstore~31 .lut_mask = 16'hCFC0;
defparam \ramstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y72_N19
dffeas \count[3] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y72_N11
dffeas \count[2] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y72_N5
dffeas \count[1] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y72_N1
dffeas \count[0] (
	.clk(\CLK~inputclkctrl_outclk ),
	.d(\count~3_combout ),
	.asdata(vcc),
	.clrn(\nRST~inputclkctrl_outclk ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N12
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// \Equal0~0_combout  = (!count[2] & (!count[3] & (!count[1] & !count[0])))

	.dataa(count[2]),
	.datab(count[3]),
	.datac(count[1]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N6
cycloneive_lcell_comb \CPUCLK~0 (
// Equation(s):
// \CPUCLK~0_combout  = \CPUCLK~q  $ (\Equal0~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\CPUCLK~q ),
	.datad(\Equal0~0_combout ),
	.cin(gnd),
	.combout(\CPUCLK~0_combout ),
	.cout());
// synopsys translate_off
defparam \CPUCLK~0 .lut_mask = 16'h0FF0;
defparam \CPUCLK~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N18
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = count[3] $ (((count[2] & (count[1] & count[0]))))

	.dataa(count[2]),
	.datab(count[1]),
	.datac(count[3]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h78F0;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N10
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = count[2] $ (((count[1] & count[0])))

	.dataa(gnd),
	.datab(count[1]),
	.datac(count[2]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h3CF0;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N4
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = count[1] $ (count[0])

	.dataa(gnd),
	.datab(gnd),
	.datac(count[1]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h0FF0;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y72_N0
cycloneive_lcell_comb \count~3 (
// Equation(s):
// \count~3_combout  = (!count[0] & ((count[2]) # ((count[1]) # (count[3]))))

	.dataa(count[2]),
	.datab(count[1]),
	.datac(count[0]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\count~3_combout ),
	.cout());
// synopsys translate_off
defparam \count~3 .lut_mask = 16'h0F0E;
defparam \count~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N4
cycloneive_lcell_comb \ramaddr~29_wirecell (
// Equation(s):
// \ramaddr~29_wirecell_combout  = !\ramaddr~29_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\ramaddr~29_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ramaddr~29_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \ramaddr~29_wirecell .lut_mask = 16'h0F0F;
defparam \ramaddr~29_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: JTAG_X1_Y37_N0
cycloneive_jtag altera_internal_jtag(
	.tms(\altera_reserved_tms~input_o ),
	.tck(\altera_reserved_tck~input_o ),
	.tdi(\altera_reserved_tdi~input_o ),
	.tdoutap(gnd),
	.tdouser(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.tdo(\altera_internal_jtag~TDO ),
	.tmsutap(\altera_internal_jtag~TMSUTAP ),
	.tckutap(\altera_internal_jtag~TCKUTAP ),
	.tdiutap(\altera_internal_jtag~TDIUTAP ),
	.shiftuser(),
	.clkdruser(),
	.updateuser(),
	.runidleuser(),
	.usr1user());

// Location: FF_X46_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y35_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y35_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y35_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y35_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X43_Y35_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .lut_mask = 16'hBB88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y35_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y35_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y35_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y35_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y35_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y35_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .lut_mask = 16'h33CC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[0]~6 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .lut_mask = 16'hC303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[1]~8 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~10 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9 .lut_mask = 16'h3CCF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[2]~10 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11 .lut_mask = 16'hA505;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y35_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[3]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13 .lut_mask = 16'h3C3C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .lut_mask = 16'hBB88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y35_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .lut_mask = 16'h55AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[0]~12 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~14 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .lut_mask = 16'hA50A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[2]~16 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18_combout ),
	.cout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .lut_mask = 16'h3C3F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[3]~19 ),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .lut_mask = 16'hA5A5;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[4]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .lut_mask = 16'hEE44;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y35_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.asdata(\altera_internal_jtag~TDIUTAP ),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .lut_mask = 16'hEE44;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y32_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y32_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y32_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y32_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y32_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0 .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y35_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .lut_mask = 16'hCC8A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .lut_mask = 16'hCC00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .lut_mask = 16'hE2AA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .lut_mask = 16'h0700;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .lut_mask = 16'hACA8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~2_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena[1]~reg0_q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .lut_mask = 16'h88D8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .lut_mask = 16'hF0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .lut_mask = 16'h0003;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .lut_mask = 16'h370C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~10_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .lut_mask = 16'hF303;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 .lut_mask = 16'h8000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .lut_mask = 16'h5F5F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .lut_mask = 16'hE0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 (
	.dataa(\altera_internal_jtag~TDIUTAP ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .lut_mask = 16'hAAF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .lut_mask = 16'hE2E2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .lut_mask = 16'hC001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~6_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .lut_mask = 16'h0010;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y35_N23
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~7_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .lut_mask = 16'hF0F8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .lut_mask = 16'h0A98;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .lut_mask = 16'hB4F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [1]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .lut_mask = 16'h4000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .lut_mask = 16'hABAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16 .lut_mask = 16'hECA0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg[4]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .lut_mask = 16'h2000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .lut_mask = 16'h0040;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .lut_mask = 16'hF546;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .lut_mask = 16'hF330;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .lut_mask = 16'hFFFE;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y35_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [2]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .lut_mask = 16'h8D88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .lut_mask = 16'h4400;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .lut_mask = 16'h0104;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y35_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg[3]~12_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .lut_mask = 16'h00F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .lut_mask = 16'hFF01;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~10_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .lut_mask = 16'h0002;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y35_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~11_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .lut_mask = 16'hAAEA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X47_Y35_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .lut_mask = 16'hB914;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~18_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .lut_mask = 16'hF5A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [2]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .lut_mask = 16'h000E;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~13_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .lut_mask = 16'h00EA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .lut_mask = 16'hFFE0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~15_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~14_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .lut_mask = 16'h434C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~17_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .lut_mask = 16'h88F8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y35_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|clear_signal~combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_dr_scan_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .lut_mask = 16'hBAAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|word_counter[1]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y35_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~9_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .lut_mask = 16'h5F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [3]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .lut_mask = 16'hA8F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|mixer_addr_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~9_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~8_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .lut_mask = 16'hF5E4;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N22
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N8
cycloneive_io_ibuf \syif.addr[1]~input (
	.i(\syif.addr [1]),
	.ibar(gnd),
	.o(\syif.addr[1]~input_o ));
// synopsys translate_off
defparam \syif.addr[1]~input .bus_hold = "false";
defparam \syif.addr[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y0_N1
cycloneive_io_ibuf \syif.tbCTRL~input (
	.i(\syif.tbCTRL ),
	.ibar(gnd),
	.o(\syif.tbCTRL~input_o ));
// synopsys translate_off
defparam \syif.tbCTRL~input .bus_hold = "false";
defparam \syif.tbCTRL~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N1
cycloneive_io_ibuf \syif.addr[0]~input (
	.i(\syif.addr [0]),
	.ibar(gnd),
	.o(\syif.addr[0]~input_o ));
// synopsys translate_off
defparam \syif.addr[0]~input .bus_hold = "false";
defparam \syif.addr[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N1
cycloneive_io_ibuf \syif.addr[3]~input (
	.i(\syif.addr [3]),
	.ibar(gnd),
	.o(\syif.addr[3]~input_o ));
// synopsys translate_off
defparam \syif.addr[3]~input .bus_hold = "false";
defparam \syif.addr[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N15
cycloneive_io_ibuf \syif.addr[2]~input (
	.i(\syif.addr [2]),
	.ibar(gnd),
	.o(\syif.addr[2]~input_o ));
// synopsys translate_off
defparam \syif.addr[2]~input .bus_hold = "false";
defparam \syif.addr[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N22
cycloneive_io_ibuf \syif.addr[5]~input (
	.i(\syif.addr [5]),
	.ibar(gnd),
	.o(\syif.addr[5]~input_o ));
// synopsys translate_off
defparam \syif.addr[5]~input .bus_hold = "false";
defparam \syif.addr[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N8
cycloneive_io_ibuf \syif.addr[4]~input (
	.i(\syif.addr [4]),
	.ibar(gnd),
	.o(\syif.addr[4]~input_o ));
// synopsys translate_off
defparam \syif.addr[4]~input .bus_hold = "false";
defparam \syif.addr[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N8
cycloneive_io_ibuf \syif.addr[7]~input (
	.i(\syif.addr [7]),
	.ibar(gnd),
	.o(\syif.addr[7]~input_o ));
// synopsys translate_off
defparam \syif.addr[7]~input .bus_hold = "false";
defparam \syif.addr[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N1
cycloneive_io_ibuf \syif.addr[6]~input (
	.i(\syif.addr [6]),
	.ibar(gnd),
	.o(\syif.addr[6]~input_o ));
// synopsys translate_off
defparam \syif.addr[6]~input .bus_hold = "false";
defparam \syif.addr[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N15
cycloneive_io_ibuf \syif.addr[9]~input (
	.i(\syif.addr [9]),
	.ibar(gnd),
	.o(\syif.addr[9]~input_o ));
// synopsys translate_off
defparam \syif.addr[9]~input .bus_hold = "false";
defparam \syif.addr[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N1
cycloneive_io_ibuf \syif.addr[8]~input (
	.i(\syif.addr [8]),
	.ibar(gnd),
	.o(\syif.addr[8]~input_o ));
// synopsys translate_off
defparam \syif.addr[8]~input .bus_hold = "false";
defparam \syif.addr[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N1
cycloneive_io_ibuf \syif.addr[11]~input (
	.i(\syif.addr [11]),
	.ibar(gnd),
	.o(\syif.addr[11]~input_o ));
// synopsys translate_off
defparam \syif.addr[11]~input .bus_hold = "false";
defparam \syif.addr[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y0_N8
cycloneive_io_ibuf \syif.addr[10]~input (
	.i(\syif.addr [10]),
	.ibar(gnd),
	.o(\syif.addr[10]~input_o ));
// synopsys translate_off
defparam \syif.addr[10]~input .bus_hold = "false";
defparam \syif.addr[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N22
cycloneive_io_ibuf \syif.addr[13]~input (
	.i(\syif.addr [13]),
	.ibar(gnd),
	.o(\syif.addr[13]~input_o ));
// synopsys translate_off
defparam \syif.addr[13]~input .bus_hold = "false";
defparam \syif.addr[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N8
cycloneive_io_ibuf \syif.addr[12]~input (
	.i(\syif.addr [12]),
	.ibar(gnd),
	.o(\syif.addr[12]~input_o ));
// synopsys translate_off
defparam \syif.addr[12]~input .bus_hold = "false";
defparam \syif.addr[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N22
cycloneive_io_ibuf \syif.addr[15]~input (
	.i(\syif.addr [15]),
	.ibar(gnd),
	.o(\syif.addr[15]~input_o ));
// synopsys translate_off
defparam \syif.addr[15]~input .bus_hold = "false";
defparam \syif.addr[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y0_N22
cycloneive_io_ibuf \syif.addr[14]~input (
	.i(\syif.addr [14]),
	.ibar(gnd),
	.o(\syif.addr[14]~input_o ));
// synopsys translate_off
defparam \syif.addr[14]~input .bus_hold = "false";
defparam \syif.addr[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N15
cycloneive_io_ibuf \syif.addr[23]~input (
	.i(\syif.addr [23]),
	.ibar(gnd),
	.o(\syif.addr[23]~input_o ));
// synopsys translate_off
defparam \syif.addr[23]~input .bus_hold = "false";
defparam \syif.addr[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N8
cycloneive_io_ibuf \syif.addr[22]~input (
	.i(\syif.addr [22]),
	.ibar(gnd),
	.o(\syif.addr[22]~input_o ));
// synopsys translate_off
defparam \syif.addr[22]~input .bus_hold = "false";
defparam \syif.addr[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N15
cycloneive_io_ibuf \syif.WEN~input (
	.i(\syif.WEN ),
	.ibar(gnd),
	.o(\syif.WEN~input_o ));
// synopsys translate_off
defparam \syif.WEN~input .bus_hold = "false";
defparam \syif.WEN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y30_N1
cycloneive_io_ibuf \syif.REN~input (
	.i(\syif.REN ),
	.ibar(gnd),
	.o(\syif.REN~input_o ));
// synopsys translate_off
defparam \syif.REN~input .bus_hold = "false";
defparam \syif.REN~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X62_Y73_N15
cycloneive_io_ibuf \syif.addr[21]~input (
	.i(\syif.addr [21]),
	.ibar(gnd),
	.o(\syif.addr[21]~input_o ));
// synopsys translate_off
defparam \syif.addr[21]~input .bus_hold = "false";
defparam \syif.addr[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y0_N22
cycloneive_io_ibuf \syif.addr[29]~input (
	.i(\syif.addr [29]),
	.ibar(gnd),
	.o(\syif.addr[29]~input_o ));
// synopsys translate_off
defparam \syif.addr[29]~input .bus_hold = "false";
defparam \syif.addr[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N22
cycloneive_io_ibuf \syif.addr[28]~input (
	.i(\syif.addr [28]),
	.ibar(gnd),
	.o(\syif.addr[28]~input_o ));
// synopsys translate_off
defparam \syif.addr[28]~input .bus_hold = "false";
defparam \syif.addr[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N1
cycloneive_io_ibuf \syif.addr[31]~input (
	.i(\syif.addr [31]),
	.ibar(gnd),
	.o(\syif.addr[31]~input_o ));
// synopsys translate_off
defparam \syif.addr[31]~input .bus_hold = "false";
defparam \syif.addr[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y29_N1
cycloneive_io_ibuf \syif.addr[30]~input (
	.i(\syif.addr [30]),
	.ibar(gnd),
	.o(\syif.addr[30]~input_o ));
// synopsys translate_off
defparam \syif.addr[30]~input .bus_hold = "false";
defparam \syif.addr[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X74_Y0_N1
cycloneive_io_ibuf \syif.addr[20]~input (
	.i(\syif.addr [20]),
	.ibar(gnd),
	.o(\syif.addr[20]~input_o ));
// synopsys translate_off
defparam \syif.addr[20]~input .bus_hold = "false";
defparam \syif.addr[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X69_Y0_N8
cycloneive_io_ibuf \syif.addr[17]~input (
	.i(\syif.addr [17]),
	.ibar(gnd),
	.o(\syif.addr[17]~input_o ));
// synopsys translate_off
defparam \syif.addr[17]~input .bus_hold = "false";
defparam \syif.addr[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y29_N8
cycloneive_io_ibuf \syif.addr[16]~input (
	.i(\syif.addr [16]),
	.ibar(gnd),
	.o(\syif.addr[16]~input_o ));
// synopsys translate_off
defparam \syif.addr[16]~input .bus_hold = "false";
defparam \syif.addr[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N15
cycloneive_io_ibuf \syif.addr[19]~input (
	.i(\syif.addr [19]),
	.ibar(gnd),
	.o(\syif.addr[19]~input_o ));
// synopsys translate_off
defparam \syif.addr[19]~input .bus_hold = "false";
defparam \syif.addr[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y29_N15
cycloneive_io_ibuf \syif.addr[18]~input (
	.i(\syif.addr [18]),
	.ibar(gnd),
	.o(\syif.addr[18]~input_o ));
// synopsys translate_off
defparam \syif.addr[18]~input .bus_hold = "false";
defparam \syif.addr[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X79_Y0_N1
cycloneive_io_ibuf \syif.addr[25]~input (
	.i(\syif.addr [25]),
	.ibar(gnd),
	.o(\syif.addr[25]~input_o ));
// synopsys translate_off
defparam \syif.addr[25]~input .bus_hold = "false";
defparam \syif.addr[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X72_Y0_N8
cycloneive_io_ibuf \syif.addr[24]~input (
	.i(\syif.addr [24]),
	.ibar(gnd),
	.o(\syif.addr[24]~input_o ));
// synopsys translate_off
defparam \syif.addr[24]~input .bus_hold = "false";
defparam \syif.addr[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X67_Y0_N1
cycloneive_io_ibuf \syif.addr[27]~input (
	.i(\syif.addr [27]),
	.ibar(gnd),
	.o(\syif.addr[27]~input_o ));
// synopsys translate_off
defparam \syif.addr[27]~input .bus_hold = "false";
defparam \syif.addr[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X60_Y73_N1
cycloneive_io_ibuf \syif.addr[26]~input (
	.i(\syif.addr [26]),
	.ibar(gnd),
	.o(\syif.addr[26]~input_o ));
// synopsys translate_off
defparam \syif.addr[26]~input .bus_hold = "false";
defparam \syif.addr[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N15
cycloneive_io_ibuf \nRST~input (
	.i(nRST),
	.ibar(gnd),
	.o(\nRST~input_o ));
// synopsys translate_off
defparam \nRST~input .bus_hold = "false";
defparam \nRST~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y36_N8
cycloneive_io_ibuf \CLK~input (
	.i(CLK),
	.ibar(gnd),
	.o(\CLK~input_o ));
// synopsys translate_off
defparam \CLK~input .bus_hold = "false";
defparam \CLK~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X33_Y0_N1
cycloneive_io_ibuf \syif.store[0]~input (
	.i(\syif.store [0]),
	.ibar(gnd),
	.o(\syif.store[0]~input_o ));
// synopsys translate_off
defparam \syif.store[0]~input .bus_hold = "false";
defparam \syif.store[0]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X47_Y73_N15
cycloneive_io_ibuf \syif.store[1]~input (
	.i(\syif.store [1]),
	.ibar(gnd),
	.o(\syif.store[1]~input_o ));
// synopsys translate_off
defparam \syif.store[1]~input .bus_hold = "false";
defparam \syif.store[1]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N22
cycloneive_io_ibuf \syif.store[2]~input (
	.i(\syif.store [2]),
	.ibar(gnd),
	.o(\syif.store[2]~input_o ));
// synopsys translate_off
defparam \syif.store[2]~input .bus_hold = "false";
defparam \syif.store[2]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N8
cycloneive_io_ibuf \syif.store[3]~input (
	.i(\syif.store [3]),
	.ibar(gnd),
	.o(\syif.store[3]~input_o ));
// synopsys translate_off
defparam \syif.store[3]~input .bus_hold = "false";
defparam \syif.store[3]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N22
cycloneive_io_ibuf \syif.store[4]~input (
	.i(\syif.store [4]),
	.ibar(gnd),
	.o(\syif.store[4]~input_o ));
// synopsys translate_off
defparam \syif.store[4]~input .bus_hold = "false";
defparam \syif.store[4]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y26_N15
cycloneive_io_ibuf \syif.store[5]~input (
	.i(\syif.store [5]),
	.ibar(gnd),
	.o(\syif.store[5]~input_o ));
// synopsys translate_off
defparam \syif.store[5]~input .bus_hold = "false";
defparam \syif.store[5]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X33_Y0_N8
cycloneive_io_ibuf \syif.store[6]~input (
	.i(\syif.store [6]),
	.ibar(gnd),
	.o(\syif.store[6]~input_o ));
// synopsys translate_off
defparam \syif.store[6]~input .bus_hold = "false";
defparam \syif.store[6]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N15
cycloneive_io_ibuf \syif.store[7]~input (
	.i(\syif.store [7]),
	.ibar(gnd),
	.o(\syif.store[7]~input_o ));
// synopsys translate_off
defparam \syif.store[7]~input .bus_hold = "false";
defparam \syif.store[7]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y0_N22
cycloneive_io_ibuf \syif.store[8]~input (
	.i(\syif.store [8]),
	.ibar(gnd),
	.o(\syif.store[8]~input_o ));
// synopsys translate_off
defparam \syif.store[8]~input .bus_hold = "false";
defparam \syif.store[8]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y29_N22
cycloneive_io_ibuf \syif.store[9]~input (
	.i(\syif.store [9]),
	.ibar(gnd),
	.o(\syif.store[9]~input_o ));
// synopsys translate_off
defparam \syif.store[9]~input .bus_hold = "false";
defparam \syif.store[9]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X42_Y0_N15
cycloneive_io_ibuf \syif.store[10]~input (
	.i(\syif.store [10]),
	.ibar(gnd),
	.o(\syif.store[10]~input_o ));
// synopsys translate_off
defparam \syif.store[10]~input .bus_hold = "false";
defparam \syif.store[10]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N1
cycloneive_io_ibuf \syif.store[11]~input (
	.i(\syif.store [11]),
	.ibar(gnd),
	.o(\syif.store[11]~input_o ));
// synopsys translate_off
defparam \syif.store[11]~input .bus_hold = "false";
defparam \syif.store[11]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y73_N22
cycloneive_io_ibuf \syif.store[12]~input (
	.i(\syif.store [12]),
	.ibar(gnd),
	.o(\syif.store[12]~input_o ));
// synopsys translate_off
defparam \syif.store[12]~input .bus_hold = "false";
defparam \syif.store[12]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X52_Y0_N15
cycloneive_io_ibuf \syif.store[13]~input (
	.i(\syif.store [13]),
	.ibar(gnd),
	.o(\syif.store[13]~input_o ));
// synopsys translate_off
defparam \syif.store[13]~input .bus_hold = "false";
defparam \syif.store[13]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y73_N15
cycloneive_io_ibuf \syif.store[14]~input (
	.i(\syif.store [14]),
	.ibar(gnd),
	.o(\syif.store[14]~input_o ));
// synopsys translate_off
defparam \syif.store[14]~input .bus_hold = "false";
defparam \syif.store[14]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y30_N1
cycloneive_io_ibuf \syif.store[15]~input (
	.i(\syif.store [15]),
	.ibar(gnd),
	.o(\syif.store[15]~input_o ));
// synopsys translate_off
defparam \syif.store[15]~input .bus_hold = "false";
defparam \syif.store[15]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y31_N15
cycloneive_io_ibuf \syif.store[16]~input (
	.i(\syif.store [16]),
	.ibar(gnd),
	.o(\syif.store[16]~input_o ));
// synopsys translate_off
defparam \syif.store[16]~input .bus_hold = "false";
defparam \syif.store[16]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y0_N15
cycloneive_io_ibuf \syif.store[17]~input (
	.i(\syif.store [17]),
	.ibar(gnd),
	.o(\syif.store[17]~input_o ));
// synopsys translate_off
defparam \syif.store[17]~input .bus_hold = "false";
defparam \syif.store[17]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X45_Y73_N8
cycloneive_io_ibuf \syif.store[18]~input (
	.i(\syif.store [18]),
	.ibar(gnd),
	.o(\syif.store[18]~input_o ));
// synopsys translate_off
defparam \syif.store[18]~input .bus_hold = "false";
defparam \syif.store[18]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X35_Y0_N22
cycloneive_io_ibuf \syif.store[19]~input (
	.i(\syif.store [19]),
	.ibar(gnd),
	.o(\syif.store[19]~input_o ));
// synopsys translate_off
defparam \syif.store[19]~input .bus_hold = "false";
defparam \syif.store[19]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N15
cycloneive_io_ibuf \syif.store[20]~input (
	.i(\syif.store [20]),
	.ibar(gnd),
	.o(\syif.store[20]~input_o ));
// synopsys translate_off
defparam \syif.store[20]~input .bus_hold = "false";
defparam \syif.store[20]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N22
cycloneive_io_ibuf \syif.store[21]~input (
	.i(\syif.store [21]),
	.ibar(gnd),
	.o(\syif.store[21]~input_o ));
// synopsys translate_off
defparam \syif.store[21]~input .bus_hold = "false";
defparam \syif.store[21]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y30_N8
cycloneive_io_ibuf \syif.store[22]~input (
	.i(\syif.store [22]),
	.ibar(gnd),
	.o(\syif.store[22]~input_o ));
// synopsys translate_off
defparam \syif.store[22]~input .bus_hold = "false";
defparam \syif.store[22]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X54_Y0_N22
cycloneive_io_ibuf \syif.store[23]~input (
	.i(\syif.store [23]),
	.ibar(gnd),
	.o(\syif.store[23]~input_o ));
// synopsys translate_off
defparam \syif.store[23]~input .bus_hold = "false";
defparam \syif.store[23]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N8
cycloneive_io_ibuf \syif.store[24]~input (
	.i(\syif.store [24]),
	.ibar(gnd),
	.o(\syif.store[24]~input_o ));
// synopsys translate_off
defparam \syif.store[24]~input .bus_hold = "false";
defparam \syif.store[24]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y30_N8
cycloneive_io_ibuf \syif.store[25]~input (
	.i(\syif.store [25]),
	.ibar(gnd),
	.o(\syif.store[25]~input_o ));
// synopsys translate_off
defparam \syif.store[25]~input .bus_hold = "false";
defparam \syif.store[25]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X49_Y0_N1
cycloneive_io_ibuf \syif.store[26]~input (
	.i(\syif.store [26]),
	.ibar(gnd),
	.o(\syif.store[26]~input_o ));
// synopsys translate_off
defparam \syif.store[26]~input .bus_hold = "false";
defparam \syif.store[26]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X58_Y73_N8
cycloneive_io_ibuf \syif.store[27]~input (
	.i(\syif.store [27]),
	.ibar(gnd),
	.o(\syif.store[27]~input_o ));
// synopsys translate_off
defparam \syif.store[27]~input .bus_hold = "false";
defparam \syif.store[27]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X65_Y73_N22
cycloneive_io_ibuf \syif.store[28]~input (
	.i(\syif.store [28]),
	.ibar(gnd),
	.o(\syif.store[28]~input_o ));
// synopsys translate_off
defparam \syif.store[28]~input .bus_hold = "false";
defparam \syif.store[28]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X35_Y0_N15
cycloneive_io_ibuf \syif.store[29]~input (
	.i(\syif.store [29]),
	.ibar(gnd),
	.o(\syif.store[29]~input_o ));
// synopsys translate_off
defparam \syif.store[29]~input .bus_hold = "false";
defparam \syif.store[29]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X115_Y28_N8
cycloneive_io_ibuf \syif.store[30]~input (
	.i(\syif.store [30]),
	.ibar(gnd),
	.o(\syif.store[30]~input_o ));
// synopsys translate_off
defparam \syif.store[30]~input .bus_hold = "false";
defparam \syif.store[30]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X40_Y0_N22
cycloneive_io_ibuf \syif.store[31]~input (
	.i(\syif.store [31]),
	.ibar(gnd),
	.o(\syif.store[31]~input_o ));
// synopsys translate_off
defparam \syif.store[31]~input .bus_hold = "false";
defparam \syif.store[31]~input .simulate_z_as = "z";
// synopsys translate_on

// Location: CLKCTRL_G4
cycloneive_clkctrl \altera_internal_jtag~TCKUTAPclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\altera_internal_jtag~TCKUTAP }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ));
// synopsys translate_off
defparam \altera_internal_jtag~TCKUTAPclkctrl .clock_type = "global clock";
defparam \altera_internal_jtag~TCKUTAPclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G13
cycloneive_clkctrl \CPUCLK~clkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CPUCLK~q }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CPUCLK~clkctrl_outclk ));
// synopsys translate_off
defparam \CPUCLK~clkctrl .clock_type = "global clock";
defparam \CPUCLK~clkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G1
cycloneive_clkctrl \nRST~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\nRST~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\nRST~inputclkctrl_outclk ));
// synopsys translate_off
defparam \nRST~inputclkctrl .clock_type = "global clock";
defparam \nRST~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: CLKCTRL_G2
cycloneive_clkctrl \CLK~inputclkctrl (
	.ena(vcc),
	.inclk({vcc,vcc,vcc,\CLK~input_o }),
	.clkselect(2'b00),
	.devclrn(devclrn),
	.devpor(devpor),
	.outclk(\CLK~inputclkctrl_outclk ));
// synopsys translate_off
defparam \CLK~inputclkctrl .clock_type = "global clock";
defparam \CLK~inputclkctrl .ena_register_mode = "none";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|node_ena_proc~1_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y35_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_shift_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|identity_contrib_update_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: IOOBUF_X38_Y0_N2
cycloneive_io_obuf \syif.halt~output (
	.i(\CPU|DP|dpif.halt~q ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.halt ),
	.obar());
// synopsys translate_off
defparam \syif.halt~output .bus_hold = "false";
defparam \syif.halt~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X49_Y0_N9
cycloneive_io_obuf \syif.load[0]~output (
	.i(\RAM|ramif.ramload[0]~0_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [0]),
	.obar());
// synopsys translate_off
defparam \syif.load[0]~output .bus_hold = "false";
defparam \syif.load[0]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y0_N2
cycloneive_io_obuf \syif.load[1]~output (
	.i(\RAM|ramif.ramload[1]~1_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [1]),
	.obar());
// synopsys translate_off
defparam \syif.load[1]~output .bus_hold = "false";
defparam \syif.load[1]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y0_N9
cycloneive_io_obuf \syif.load[2]~output (
	.i(\RAM|ramif.ramload[2]~2_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [2]),
	.obar());
// synopsys translate_off
defparam \syif.load[2]~output .bus_hold = "false";
defparam \syif.load[2]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X38_Y0_N9
cycloneive_io_obuf \syif.load[3]~output (
	.i(\RAM|ramif.ramload[3]~3_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [3]),
	.obar());
// synopsys translate_off
defparam \syif.load[3]~output .bus_hold = "false";
defparam \syif.load[3]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y27_N16
cycloneive_io_obuf \syif.load[4]~output (
	.i(\RAM|ramif.ramload[4]~4_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [4]),
	.obar());
// synopsys translate_off
defparam \syif.load[4]~output .bus_hold = "false";
defparam \syif.load[4]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X79_Y0_N23
cycloneive_io_obuf \syif.load[5]~output (
	.i(\RAM|ramif.ramload[5]~5_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [5]),
	.obar());
// synopsys translate_off
defparam \syif.load[5]~output .bus_hold = "false";
defparam \syif.load[5]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y28_N23
cycloneive_io_obuf \syif.load[6]~output (
	.i(\RAM|ramif.ramload[6]~6_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [6]),
	.obar());
// synopsys translate_off
defparam \syif.load[6]~output .bus_hold = "false";
defparam \syif.load[6]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N16
cycloneive_io_obuf \syif.load[7]~output (
	.i(\RAM|ramif.ramload[7]~7_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [7]),
	.obar());
// synopsys translate_off
defparam \syif.load[7]~output .bus_hold = "false";
defparam \syif.load[7]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X79_Y0_N9
cycloneive_io_obuf \syif.load[8]~output (
	.i(\RAM|ramif.ramload[8]~8_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [8]),
	.obar());
// synopsys translate_off
defparam \syif.load[8]~output .bus_hold = "false";
defparam \syif.load[8]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y28_N2
cycloneive_io_obuf \syif.load[9]~output (
	.i(\RAM|ramif.ramload[9]~9_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [9]),
	.obar());
// synopsys translate_off
defparam \syif.load[9]~output .bus_hold = "false";
defparam \syif.load[9]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N9
cycloneive_io_obuf \syif.load[10]~output (
	.i(\RAM|ramif.ramload[10]~10_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [10]),
	.obar());
// synopsys translate_off
defparam \syif.load[10]~output .bus_hold = "false";
defparam \syif.load[10]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N16
cycloneive_io_obuf \syif.load[11]~output (
	.i(\RAM|ramif.ramload[11]~11_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [11]),
	.obar());
// synopsys translate_off
defparam \syif.load[11]~output .bus_hold = "false";
defparam \syif.load[11]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N23
cycloneive_io_obuf \syif.load[12]~output (
	.i(\RAM|ramif.ramload[12]~12_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [12]),
	.obar());
// synopsys translate_off
defparam \syif.load[12]~output .bus_hold = "false";
defparam \syif.load[12]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X52_Y73_N2
cycloneive_io_obuf \syif.load[13]~output (
	.i(\RAM|ramif.ramload[13]~13_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [13]),
	.obar());
// synopsys translate_off
defparam \syif.load[13]~output .bus_hold = "false";
defparam \syif.load[13]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N9
cycloneive_io_obuf \syif.load[14]~output (
	.i(\RAM|ramif.ramload[14]~14_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [14]),
	.obar());
// synopsys translate_off
defparam \syif.load[14]~output .bus_hold = "false";
defparam \syif.load[14]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y32_N23
cycloneive_io_obuf \syif.load[15]~output (
	.i(\RAM|ramif.ramload[15]~15_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [15]),
	.obar());
// synopsys translate_off
defparam \syif.load[15]~output .bus_hold = "false";
defparam \syif.load[15]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X67_Y0_N16
cycloneive_io_obuf \syif.load[16]~output (
	.i(\RAM|ramif.ramload[16]~16_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [16]),
	.obar());
// synopsys translate_off
defparam \syif.load[16]~output .bus_hold = "false";
defparam \syif.load[16]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y73_N9
cycloneive_io_obuf \syif.load[17]~output (
	.i(\RAM|ramif.ramload[17]~17_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [17]),
	.obar());
// synopsys translate_off
defparam \syif.load[17]~output .bus_hold = "false";
defparam \syif.load[17]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N2
cycloneive_io_obuf \syif.load[18]~output (
	.i(\RAM|ramif.ramload[18]~18_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [18]),
	.obar());
// synopsys translate_off
defparam \syif.load[18]~output .bus_hold = "false";
defparam \syif.load[18]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X54_Y73_N9
cycloneive_io_obuf \syif.load[19]~output (
	.i(\RAM|ramif.ramload[19]~19_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [19]),
	.obar());
// synopsys translate_off
defparam \syif.load[19]~output .bus_hold = "false";
defparam \syif.load[19]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X47_Y73_N2
cycloneive_io_obuf \syif.load[20]~output (
	.i(\RAM|ramif.ramload[20]~20_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [20]),
	.obar());
// synopsys translate_off
defparam \syif.load[20]~output .bus_hold = "false";
defparam \syif.load[20]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X65_Y0_N16
cycloneive_io_obuf \syif.load[21]~output (
	.i(\RAM|ramif.ramload[21]~21_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [21]),
	.obar());
// synopsys translate_off
defparam \syif.load[21]~output .bus_hold = "false";
defparam \syif.load[21]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y73_N23
cycloneive_io_obuf \syif.load[22]~output (
	.i(\RAM|ramif.ramload[22]~22_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [22]),
	.obar());
// synopsys translate_off
defparam \syif.load[22]~output .bus_hold = "false";
defparam \syif.load[22]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X62_Y0_N16
cycloneive_io_obuf \syif.load[23]~output (
	.i(\RAM|ramif.ramload[23]~23_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [23]),
	.obar());
// synopsys translate_off
defparam \syif.load[23]~output .bus_hold = "false";
defparam \syif.load[23]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X60_Y0_N23
cycloneive_io_obuf \syif.load[24]~output (
	.i(\RAM|ramif.ramload[24]~24_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [24]),
	.obar());
// synopsys translate_off
defparam \syif.load[24]~output .bus_hold = "false";
defparam \syif.load[24]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y28_N16
cycloneive_io_obuf \syif.load[25]~output (
	.i(\RAM|ramif.ramload[25]~25_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [25]),
	.obar());
// synopsys translate_off
defparam \syif.load[25]~output .bus_hold = "false";
defparam \syif.load[25]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y27_N23
cycloneive_io_obuf \syif.load[26]~output (
	.i(\RAM|ramif.ramload[26]~26_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [26]),
	.obar());
// synopsys translate_off
defparam \syif.load[26]~output .bus_hold = "false";
defparam \syif.load[26]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N2
cycloneive_io_obuf \syif.load[27]~output (
	.i(\RAM|ramif.ramload[27]~27_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [27]),
	.obar());
// synopsys translate_off
defparam \syif.load[27]~output .bus_hold = "false";
defparam \syif.load[27]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X81_Y0_N16
cycloneive_io_obuf \syif.load[28]~output (
	.i(\RAM|ramif.ramload[28]~28_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [28]),
	.obar());
// synopsys translate_off
defparam \syif.load[28]~output .bus_hold = "false";
defparam \syif.load[28]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X56_Y0_N23
cycloneive_io_obuf \syif.load[29]~output (
	.i(\RAM|ramif.ramload[29]~29_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [29]),
	.obar());
// synopsys translate_off
defparam \syif.load[29]~output .bus_hold = "false";
defparam \syif.load[29]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X79_Y0_N16
cycloneive_io_obuf \syif.load[30]~output (
	.i(\RAM|ramif.ramload[30]~30_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [30]),
	.obar());
// synopsys translate_off
defparam \syif.load[30]~output .bus_hold = "false";
defparam \syif.load[30]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X115_Y31_N2
cycloneive_io_obuf \syif.load[31]~output (
	.i(\RAM|ramif.ramload[31]~31_combout ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(\syif.load [31]),
	.obar());
// synopsys translate_off
defparam \syif.load[31]~output .bus_hold = "false";
defparam \syif.load[31]~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOOBUF_X0_Y37_N1
cycloneive_io_obuf \altera_reserved_tdo~output (
	.i(\altera_internal_jtag~TDO ),
	.oe(vcc),
	.seriesterminationcontrol(16'b0000000000000000),
	.devoe(devoe),
	.o(altera_reserved_tdo),
	.obar());
// synopsys translate_off
defparam \altera_reserved_tdo~output .bus_hold = "false";
defparam \altera_reserved_tdo~output .open_drain_output = "false";
// synopsys translate_on

// Location: IOIBUF_X0_Y38_N1
cycloneive_io_ibuf \altera_reserved_tms~input (
	.i(altera_reserved_tms),
	.ibar(gnd),
	.o(\altera_reserved_tms~input_o ));
// synopsys translate_off
defparam \altera_reserved_tms~input .bus_hold = "false";
defparam \altera_reserved_tms~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y39_N1
cycloneive_io_ibuf \altera_reserved_tck~input (
	.i(altera_reserved_tck),
	.ibar(gnd),
	.o(\altera_reserved_tck~input_o ));
// synopsys translate_off
defparam \altera_reserved_tck~input .bus_hold = "false";
defparam \altera_reserved_tck~input .simulate_z_as = "z";
// synopsys translate_on

// Location: IOIBUF_X0_Y40_N1
cycloneive_io_ibuf \altera_reserved_tdi~input (
	.i(altera_reserved_tdi),
	.ibar(gnd),
	.o(\altera_reserved_tdi~input_o ));
// synopsys translate_off
defparam \altera_reserved_tdi~input .bus_hold = "false";
defparam \altera_reserved_tdi~input .simulate_z_as = "z";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\altera_internal_jtag~TDIUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datad(\altera_internal_jtag~TMSUTAP ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .lut_mask = 16'h0F00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .lut_mask = 16'h0FF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X49_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .lut_mask = 16'h3CF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X49_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(!\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [9]),
	.datab(\altera_internal_jtag~TMSUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|tms_cnt [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .lut_mask = 16'h3373;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .lut_mask = 16'hF0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N25
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .lut_mask = 16'hFFF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [13]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .lut_mask = 16'hC0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [10]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .lut_mask = 16'hFFFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X45_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N7
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .lut_mask = 16'hFF00;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3]~feeder_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2]~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [4]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .lut_mask = 16'h0004;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(gnd),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [2]),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [11]),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [8]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [9]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [6]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .lut_mask = 16'h0001;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|jtag_ir_reg [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal0~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .lut_mask = 16'h0400;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N20
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [14]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [12]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .lut_mask = 16'hE0E0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal1~0_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [2]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .lut_mask = 16'h0A0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .lut_mask = 16'hFA0A;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [6]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .lut_mask = 16'hA0A0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .lut_mask = 16'hFFFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y34_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .lut_mask = 16'hA080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 (
	.dataa(gnd),
	.datab(\altera_internal_jtag~TDIUTAP ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .lut_mask = 16'hCCF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N4
cycloneive_lcell_comb \~QIC_CREATED_GND~I (
// Equation(s):
// \~QIC_CREATED_GND~I_combout  = GND

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\~QIC_CREATED_GND~I_combout ),
	.cout());
// synopsys translate_off
defparam \~QIC_CREATED_GND~I .lut_mask = 16'h0000;
defparam \~QIC_CREATED_GND~I .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5]~0_combout ),
	.asdata(\~QIC_CREATED_GND~I_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N14
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~2_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg~q ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .lut_mask = 16'h30B8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N15
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2]~3_combout ),
	.asdata(vcc),
	.clrn(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y33_N21
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_dr_scan_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [7]),
	.datac(\altera_internal_jtag~TMSUTAP ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .lut_mask = 16'hF0C0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N5
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [15]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .lut_mask = 16'hFFFD;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\altera_internal_jtag~TMSUTAP ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y33_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .lut_mask = 16'hF000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y33_N1
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg_proc~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .lut_mask = 16'hB080;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y32_N17
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~6_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N30
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|is_in_use_reg~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .lut_mask = 16'hFC0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y32_N31
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~2_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N16
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~3_combout ),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .lut_mask = 16'hFAF0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N6
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 (
	.dataa(\RAM|altsyncram_component|auto_generated|mgl_prim2|tdo~1_combout ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .lut_mask = 16'hAACC;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N0
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .lut_mask = 16'h5000;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|Equal3~0_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|reset_ena_reg_proc~0_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .lut_mask = 16'h44F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N19
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0]~4_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_mode_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .lut_mask = 16'h00F0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y33_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2]~3_combout ),
	.datab(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [2]),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~7_combout ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .lut_mask = 16'hDD88;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 (
	.dataa(gnd),
	.datab(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .lut_mask = 16'hCFC0;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y32_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~9_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N18
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [4]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .lut_mask = 16'hFC0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y33_N9
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3]~1_combout ),
	.asdata(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~8_combout ),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|virtual_ir_scan_reg~q ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 (
	.dataa(gnd),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [3]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datad(\RAM|altsyncram_component|auto_generated|mgl_prim2|ir_loaded_address_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .lut_mask = 16'hFC0C;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y32_N27
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[0]~4_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y34_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\altera_internal_jtag~TDIUTAP ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .lut_mask = 16'h5050;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N24
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [4]),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .lut_mask = 16'hFAFA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X47_Y34_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N12
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [3]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .lut_mask = 16'hFFAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y34_N13
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [2]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .lut_mask = 16'h5500;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y34_N3
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y34_N10
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [3]),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [1]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .lut_mask = 16'hFFAA;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y34_N11
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] (
	.clk(\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N26
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg|WORD_SR [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [2]),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_minor_ver_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .lut_mask = 16'hF2C2;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo_bypass_reg~q ),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~1_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~0_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [5]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .lut_mask = 16'hCCB8;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y35_N28
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 (
	.dataa(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|design_hash_reg [0]),
	.datab(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~4_combout ),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~2_combout ),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irsr_reg [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .lut_mask = 16'h13CF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y35_N29
dffeas \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo (
	.clk(!\altera_internal_jtag~TCKUTAPclkctrl_outclk ),
	.d(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~5_combout ),
	.asdata(vcc),
	.clrn(!\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [8]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|hub_info_reg_ena~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.prn(vcc));
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .is_wysiwyg = "true";
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X17_Y35_N8
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~q ),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|tdo~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X1_Y63_N0
cycloneive_lcell_comb \auto_hub|~GND (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|~GND~combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|~GND .lut_mask = 16'h0000;
defparam \auto_hub|~GND .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N2
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~q ),
	.datad(gnd),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .lut_mask = 16'h0F0F;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|clr_reg~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y33_N4
cycloneive_lcell_comb \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [0]),
	.cin(gnd),
	.combout(\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell_combout ),
	.cout());
// synopsys translate_off
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .lut_mask = 16'h00FF;
defparam \auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state[0]~_wirecell .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline (
	prifdmemaddr_1,
	pc_1,
	prifdmemren,
	prifdmemwen,
	prifdmemaddr_0,
	pc_0,
	prifdmemaddr_3,
	prifdmemaddr_2,
	prifdmemaddr_5,
	prifdmemaddr_4,
	prifdmemaddr_7,
	prifdmemaddr_6,
	prifdmemaddr_9,
	prifdmemaddr_8,
	prifdmemaddr_11,
	prifdmemaddr_10,
	prifdmemaddr_13,
	prifdmemaddr_12,
	prifdmemaddr_15,
	prifdmemaddr_14,
	prifdmemaddr_23,
	prifdmemaddr_22,
	prifdmemaddr_21,
	prifdmemaddr_29,
	prifdmemaddr_28,
	prifdmemaddr_31,
	prifdmemaddr_30,
	prifdmemaddr_20,
	prifdmemaddr_17,
	prifdmemaddr_16,
	prifdmemaddr_19,
	prifdmemaddr_18,
	prifdmemaddr_25,
	prifdmemaddr_24,
	prifdmemaddr_27,
	prifdmemaddr_26,
	prifdmemstore_0,
	prifdmemstore_1,
	prifdmemstore_2,
	prifdmemstore_3,
	prifdmemstore_4,
	prifdmemstore_5,
	prifdmemstore_6,
	prifdmemstore_7,
	prifdmemstore_8,
	prifdmemstore_9,
	prifdmemstore_10,
	prifdmemstore_11,
	prifdmemstore_12,
	prifdmemstore_13,
	prifdmemstore_14,
	prifdmemstore_15,
	prifdmemstore_16,
	prifdmemstore_17,
	prifdmemstore_18,
	prifdmemstore_19,
	prifdmemstore_20,
	prifdmemstore_21,
	prifdmemstore_22,
	prifdmemstore_23,
	prifdmemstore_24,
	prifdmemstore_25,
	prifdmemstore_26,
	prifdmemstore_27,
	prifdmemstore_28,
	prifdmemstore_29,
	prifdmemstore_30,
	prifdmemstore_31,
	LessThan1,
	pc_3,
	pc_2,
	pc_5,
	pc_4,
	pc_7,
	pc_6,
	pc_9,
	pc_8,
	pc_11,
	pc_10,
	pc_13,
	pc_12,
	pc_15,
	pc_14,
	pc_23,
	pc_22,
	pc_21,
	pc_29,
	pc_28,
	pc_31,
	pc_30,
	pc_20,
	pc_17,
	pc_16,
	pc_19,
	pc_18,
	pc_25,
	pc_24,
	pc_27,
	pc_26,
	always0,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	nRST,
	CLK,
	nRST1,
	dpifhalt,
	devpor,
	devclrn,
	devoe);
output 	prifdmemaddr_1;
output 	pc_1;
output 	prifdmemren;
output 	prifdmemwen;
output 	prifdmemaddr_0;
output 	pc_0;
output 	prifdmemaddr_3;
output 	prifdmemaddr_2;
output 	prifdmemaddr_5;
output 	prifdmemaddr_4;
output 	prifdmemaddr_7;
output 	prifdmemaddr_6;
output 	prifdmemaddr_9;
output 	prifdmemaddr_8;
output 	prifdmemaddr_11;
output 	prifdmemaddr_10;
output 	prifdmemaddr_13;
output 	prifdmemaddr_12;
output 	prifdmemaddr_15;
output 	prifdmemaddr_14;
output 	prifdmemaddr_23;
output 	prifdmemaddr_22;
output 	prifdmemaddr_21;
output 	prifdmemaddr_29;
output 	prifdmemaddr_28;
output 	prifdmemaddr_31;
output 	prifdmemaddr_30;
output 	prifdmemaddr_20;
output 	prifdmemaddr_17;
output 	prifdmemaddr_16;
output 	prifdmemaddr_19;
output 	prifdmemaddr_18;
output 	prifdmemaddr_25;
output 	prifdmemaddr_24;
output 	prifdmemaddr_27;
output 	prifdmemaddr_26;
output 	prifdmemstore_0;
output 	prifdmemstore_1;
output 	prifdmemstore_2;
output 	prifdmemstore_3;
output 	prifdmemstore_4;
output 	prifdmemstore_5;
output 	prifdmemstore_6;
output 	prifdmemstore_7;
output 	prifdmemstore_8;
output 	prifdmemstore_9;
output 	prifdmemstore_10;
output 	prifdmemstore_11;
output 	prifdmemstore_12;
output 	prifdmemstore_13;
output 	prifdmemstore_14;
output 	prifdmemstore_15;
output 	prifdmemstore_16;
output 	prifdmemstore_17;
output 	prifdmemstore_18;
output 	prifdmemstore_19;
output 	prifdmemstore_20;
output 	prifdmemstore_21;
output 	prifdmemstore_22;
output 	prifdmemstore_23;
output 	prifdmemstore_24;
output 	prifdmemstore_25;
output 	prifdmemstore_26;
output 	prifdmemstore_27;
output 	prifdmemstore_28;
output 	prifdmemstore_29;
output 	prifdmemstore_30;
output 	prifdmemstore_31;
input 	LessThan1;
output 	pc_3;
output 	pc_2;
output 	pc_5;
output 	pc_4;
output 	pc_7;
output 	pc_6;
output 	pc_9;
output 	pc_8;
output 	pc_11;
output 	pc_10;
output 	pc_13;
output 	pc_12;
output 	pc_15;
output 	pc_14;
output 	pc_23;
output 	pc_22;
output 	pc_21;
output 	pc_29;
output 	pc_28;
output 	pc_31;
output 	pc_30;
output 	pc_20;
output 	pc_17;
output 	pc_16;
output 	pc_19;
output 	pc_18;
output 	pc_25;
output 	pc_24;
output 	pc_27;
output 	pc_26;
input 	always0;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	nRST;
input 	CLK;
input 	nRST1;
output 	dpifhalt;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \CC|always0~0_combout ;
wire \CC|ccif.iwait[0]~0_combout ;


memory_control CC(
	.prifdmemren(prifdmemren),
	.prifdmemwen(prifdmemwen),
	.LessThan1(LessThan1),
	.always0(always0),
	.always01(\CC|always0~0_combout ),
	.ccifiwait_0(\CC|ccif.iwait[0]~0_combout ),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

datapath DP(
	.prifdmemaddr_1(prifdmemaddr_1),
	.pc_1(pc_1),
	.prifdmemren(prifdmemren),
	.prifdmemwen(prifdmemwen),
	.prifdmemaddr_0(prifdmemaddr_0),
	.pc_0(pc_0),
	.prifdmemaddr_3(prifdmemaddr_3),
	.prifdmemaddr_2(prifdmemaddr_2),
	.prifdmemaddr_5(prifdmemaddr_5),
	.prifdmemaddr_4(prifdmemaddr_4),
	.prifdmemaddr_7(prifdmemaddr_7),
	.prifdmemaddr_6(prifdmemaddr_6),
	.prifdmemaddr_9(prifdmemaddr_9),
	.prifdmemaddr_8(prifdmemaddr_8),
	.prifdmemaddr_11(prifdmemaddr_11),
	.prifdmemaddr_10(prifdmemaddr_10),
	.prifdmemaddr_13(prifdmemaddr_13),
	.prifdmemaddr_12(prifdmemaddr_12),
	.prifdmemaddr_15(prifdmemaddr_15),
	.prifdmemaddr_14(prifdmemaddr_14),
	.prifdmemaddr_23(prifdmemaddr_23),
	.prifdmemaddr_22(prifdmemaddr_22),
	.prifdmemaddr_21(prifdmemaddr_21),
	.prifdmemaddr_29(prifdmemaddr_29),
	.prifdmemaddr_28(prifdmemaddr_28),
	.prifdmemaddr_31(prifdmemaddr_31),
	.prifdmemaddr_30(prifdmemaddr_30),
	.prifdmemaddr_20(prifdmemaddr_20),
	.prifdmemaddr_17(prifdmemaddr_17),
	.prifdmemaddr_16(prifdmemaddr_16),
	.prifdmemaddr_19(prifdmemaddr_19),
	.prifdmemaddr_18(prifdmemaddr_18),
	.prifdmemaddr_25(prifdmemaddr_25),
	.prifdmemaddr_24(prifdmemaddr_24),
	.prifdmemaddr_27(prifdmemaddr_27),
	.prifdmemaddr_26(prifdmemaddr_26),
	.prifdmemstore_0(prifdmemstore_0),
	.prifdmemstore_1(prifdmemstore_1),
	.prifdmemstore_2(prifdmemstore_2),
	.prifdmemstore_3(prifdmemstore_3),
	.prifdmemstore_4(prifdmemstore_4),
	.prifdmemstore_5(prifdmemstore_5),
	.prifdmemstore_6(prifdmemstore_6),
	.prifdmemstore_7(prifdmemstore_7),
	.prifdmemstore_8(prifdmemstore_8),
	.prifdmemstore_9(prifdmemstore_9),
	.prifdmemstore_10(prifdmemstore_10),
	.prifdmemstore_11(prifdmemstore_11),
	.prifdmemstore_12(prifdmemstore_12),
	.prifdmemstore_13(prifdmemstore_13),
	.prifdmemstore_14(prifdmemstore_14),
	.prifdmemstore_15(prifdmemstore_15),
	.prifdmemstore_16(prifdmemstore_16),
	.prifdmemstore_17(prifdmemstore_17),
	.prifdmemstore_18(prifdmemstore_18),
	.prifdmemstore_19(prifdmemstore_19),
	.prifdmemstore_20(prifdmemstore_20),
	.prifdmemstore_21(prifdmemstore_21),
	.prifdmemstore_22(prifdmemstore_22),
	.prifdmemstore_23(prifdmemstore_23),
	.prifdmemstore_24(prifdmemstore_24),
	.prifdmemstore_25(prifdmemstore_25),
	.prifdmemstore_26(prifdmemstore_26),
	.prifdmemstore_27(prifdmemstore_27),
	.prifdmemstore_28(prifdmemstore_28),
	.prifdmemstore_29(prifdmemstore_29),
	.prifdmemstore_30(prifdmemstore_30),
	.prifdmemstore_31(prifdmemstore_31),
	.LessThan1(LessThan1),
	.pc_3(pc_3),
	.pc_2(pc_2),
	.pc_5(pc_5),
	.pc_4(pc_4),
	.pc_7(pc_7),
	.pc_6(pc_6),
	.pc_9(pc_9),
	.pc_8(pc_8),
	.pc_11(pc_11),
	.pc_10(pc_10),
	.pc_13(pc_13),
	.pc_12(pc_12),
	.pc_15(pc_15),
	.pc_14(pc_14),
	.pc_23(pc_23),
	.pc_22(pc_22),
	.pc_21(pc_21),
	.pc_29(pc_29),
	.pc_28(pc_28),
	.pc_31(pc_31),
	.pc_30(pc_30),
	.pc_20(pc_20),
	.pc_17(pc_17),
	.pc_16(pc_16),
	.pc_19(pc_19),
	.pc_18(pc_18),
	.pc_25(pc_25),
	.pc_24(pc_24),
	.pc_27(pc_27),
	.pc_26(pc_26),
	.always0(always0),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.always01(\CC|always0~0_combout ),
	.ccifiwait_0(\CC|ccif.iwait[0]~0_combout ),
	.nRST(nRST),
	.CLK(CLK),
	.nRST1(nRST1),
	.dpifhalt(dpifhalt),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module datapath (
	prifdmemaddr_1,
	pc_1,
	prifdmemren,
	prifdmemwen,
	prifdmemaddr_0,
	pc_0,
	prifdmemaddr_3,
	prifdmemaddr_2,
	prifdmemaddr_5,
	prifdmemaddr_4,
	prifdmemaddr_7,
	prifdmemaddr_6,
	prifdmemaddr_9,
	prifdmemaddr_8,
	prifdmemaddr_11,
	prifdmemaddr_10,
	prifdmemaddr_13,
	prifdmemaddr_12,
	prifdmemaddr_15,
	prifdmemaddr_14,
	prifdmemaddr_23,
	prifdmemaddr_22,
	prifdmemaddr_21,
	prifdmemaddr_29,
	prifdmemaddr_28,
	prifdmemaddr_31,
	prifdmemaddr_30,
	prifdmemaddr_20,
	prifdmemaddr_17,
	prifdmemaddr_16,
	prifdmemaddr_19,
	prifdmemaddr_18,
	prifdmemaddr_25,
	prifdmemaddr_24,
	prifdmemaddr_27,
	prifdmemaddr_26,
	prifdmemstore_0,
	prifdmemstore_1,
	prifdmemstore_2,
	prifdmemstore_3,
	prifdmemstore_4,
	prifdmemstore_5,
	prifdmemstore_6,
	prifdmemstore_7,
	prifdmemstore_8,
	prifdmemstore_9,
	prifdmemstore_10,
	prifdmemstore_11,
	prifdmemstore_12,
	prifdmemstore_13,
	prifdmemstore_14,
	prifdmemstore_15,
	prifdmemstore_16,
	prifdmemstore_17,
	prifdmemstore_18,
	prifdmemstore_19,
	prifdmemstore_20,
	prifdmemstore_21,
	prifdmemstore_22,
	prifdmemstore_23,
	prifdmemstore_24,
	prifdmemstore_25,
	prifdmemstore_26,
	prifdmemstore_27,
	prifdmemstore_28,
	prifdmemstore_29,
	prifdmemstore_30,
	prifdmemstore_31,
	LessThan1,
	pc_3,
	pc_2,
	pc_5,
	pc_4,
	pc_7,
	pc_6,
	pc_9,
	pc_8,
	pc_11,
	pc_10,
	pc_13,
	pc_12,
	pc_15,
	pc_14,
	pc_23,
	pc_22,
	pc_21,
	pc_29,
	pc_28,
	pc_31,
	pc_30,
	pc_20,
	pc_17,
	pc_16,
	pc_19,
	pc_18,
	pc_25,
	pc_24,
	pc_27,
	pc_26,
	always0,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	always01,
	ccifiwait_0,
	nRST,
	CLK,
	nRST1,
	dpifhalt,
	devpor,
	devclrn,
	devoe);
output 	prifdmemaddr_1;
output 	pc_1;
output 	prifdmemren;
output 	prifdmemwen;
output 	prifdmemaddr_0;
output 	pc_0;
output 	prifdmemaddr_3;
output 	prifdmemaddr_2;
output 	prifdmemaddr_5;
output 	prifdmemaddr_4;
output 	prifdmemaddr_7;
output 	prifdmemaddr_6;
output 	prifdmemaddr_9;
output 	prifdmemaddr_8;
output 	prifdmemaddr_11;
output 	prifdmemaddr_10;
output 	prifdmemaddr_13;
output 	prifdmemaddr_12;
output 	prifdmemaddr_15;
output 	prifdmemaddr_14;
output 	prifdmemaddr_23;
output 	prifdmemaddr_22;
output 	prifdmemaddr_21;
output 	prifdmemaddr_29;
output 	prifdmemaddr_28;
output 	prifdmemaddr_31;
output 	prifdmemaddr_30;
output 	prifdmemaddr_20;
output 	prifdmemaddr_17;
output 	prifdmemaddr_16;
output 	prifdmemaddr_19;
output 	prifdmemaddr_18;
output 	prifdmemaddr_25;
output 	prifdmemaddr_24;
output 	prifdmemaddr_27;
output 	prifdmemaddr_26;
output 	prifdmemstore_0;
output 	prifdmemstore_1;
output 	prifdmemstore_2;
output 	prifdmemstore_3;
output 	prifdmemstore_4;
output 	prifdmemstore_5;
output 	prifdmemstore_6;
output 	prifdmemstore_7;
output 	prifdmemstore_8;
output 	prifdmemstore_9;
output 	prifdmemstore_10;
output 	prifdmemstore_11;
output 	prifdmemstore_12;
output 	prifdmemstore_13;
output 	prifdmemstore_14;
output 	prifdmemstore_15;
output 	prifdmemstore_16;
output 	prifdmemstore_17;
output 	prifdmemstore_18;
output 	prifdmemstore_19;
output 	prifdmemstore_20;
output 	prifdmemstore_21;
output 	prifdmemstore_22;
output 	prifdmemstore_23;
output 	prifdmemstore_24;
output 	prifdmemstore_25;
output 	prifdmemstore_26;
output 	prifdmemstore_27;
output 	prifdmemstore_28;
output 	prifdmemstore_29;
output 	prifdmemstore_30;
output 	prifdmemstore_31;
input 	LessThan1;
output 	pc_3;
output 	pc_2;
output 	pc_5;
output 	pc_4;
output 	pc_7;
output 	pc_6;
output 	pc_9;
output 	pc_8;
output 	pc_11;
output 	pc_10;
output 	pc_13;
output 	pc_12;
output 	pc_15;
output 	pc_14;
output 	pc_23;
output 	pc_22;
output 	pc_21;
output 	pc_29;
output 	pc_28;
output 	pc_31;
output 	pc_30;
output 	pc_20;
output 	pc_17;
output 	pc_16;
output 	pc_19;
output 	pc_18;
output 	pc_25;
output 	pc_24;
output 	pc_27;
output 	pc_26;
input 	always0;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	always01;
input 	ccifiwait_0;
input 	nRST;
input 	CLK;
input 	nRST1;
output 	dpifhalt;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \prif.Regwen_mem~q ;
wire \prif.memren_ex~q ;
wire \prif.memwen_ex~q ;
wire \Add3~14_combout ;
wire \Add3~30_combout ;
wire \Add3~34_combout ;
wire \Add3~46_combout ;
wire \prif.halt_ex~q ;
wire \prif.Regwen_ex~q ;
wire \Add0~1 ;
wire \Add0~0_combout ;
wire \Add0~3 ;
wire \Add0~2_combout ;
wire \Add0~5 ;
wire \Add0~4_combout ;
wire \Add0~7 ;
wire \Add0~6_combout ;
wire \Add0~9 ;
wire \Add0~8_combout ;
wire \Add0~11 ;
wire \Add0~10_combout ;
wire \Add0~13 ;
wire \Add0~12_combout ;
wire \Add0~15 ;
wire \Add0~14_combout ;
wire \Add0~17 ;
wire \Add0~16_combout ;
wire \Add0~19 ;
wire \Add0~18_combout ;
wire \Add0~21 ;
wire \Add0~20_combout ;
wire \Add0~23 ;
wire \Add0~22_combout ;
wire \Add0~25 ;
wire \Add0~24_combout ;
wire \Add0~27 ;
wire \Add0~26_combout ;
wire \Add0~29 ;
wire \Add0~28_combout ;
wire \Add0~31 ;
wire \Add0~30_combout ;
wire \Add0~33 ;
wire \Add0~32_combout ;
wire \Add0~35 ;
wire \Add0~34_combout ;
wire \Add0~37 ;
wire \Add0~36_combout ;
wire \Add0~39 ;
wire \Add0~38_combout ;
wire \Add0~41 ;
wire \Add0~40_combout ;
wire \Add0~43 ;
wire \Add0~42_combout ;
wire \Add0~45 ;
wire \Add0~44_combout ;
wire \Add0~47 ;
wire \Add0~46_combout ;
wire \Add0~49 ;
wire \Add0~48_combout ;
wire \Add0~51 ;
wire \Add0~50_combout ;
wire \Add0~53 ;
wire \Add0~52_combout ;
wire \Add0~55 ;
wire \Add0~54_combout ;
wire \Add0~57 ;
wire \Add0~56_combout ;
wire \Add0~58_combout ;
wire \Add2~1 ;
wire \Add2~0_combout ;
wire \Add2~3 ;
wire \Add2~2_combout ;
wire \Add2~5 ;
wire \Add2~4_combout ;
wire \Add2~7 ;
wire \Add2~6_combout ;
wire \Add2~9 ;
wire \Add2~8_combout ;
wire \Add2~11 ;
wire \Add2~10_combout ;
wire \Add2~13 ;
wire \Add2~12_combout ;
wire \Add2~15 ;
wire \Add2~14_combout ;
wire \Add2~17 ;
wire \Add2~16_combout ;
wire \Add2~19 ;
wire \Add2~18_combout ;
wire \Add2~21 ;
wire \Add2~20_combout ;
wire \Add2~23 ;
wire \Add2~22_combout ;
wire \Add2~25 ;
wire \Add2~24_combout ;
wire \Add2~27 ;
wire \Add2~26_combout ;
wire \Add2~29 ;
wire \Add2~28_combout ;
wire \Add2~31 ;
wire \Add2~30_combout ;
wire \Add2~33 ;
wire \Add2~32_combout ;
wire \Add2~35 ;
wire \Add2~34_combout ;
wire \Add2~37 ;
wire \Add2~36_combout ;
wire \Add2~39 ;
wire \Add2~38_combout ;
wire \Add2~41 ;
wire \Add2~40_combout ;
wire \Add2~43 ;
wire \Add2~42_combout ;
wire \Add2~45 ;
wire \Add2~44_combout ;
wire \Add2~47 ;
wire \Add2~46_combout ;
wire \Add2~49 ;
wire \Add2~48_combout ;
wire \Add2~51 ;
wire \Add2~50_combout ;
wire \Add2~53 ;
wire \Add2~52_combout ;
wire \Add2~55 ;
wire \Add2~54_combout ;
wire \Add2~56_combout ;
wire \Mux94~0_combout ;
wire \Mux89~2_combout ;
wire \HU|ptBScr~1_combout ;
wire \prif.Regwen_wb~q ;
wire \HU|Equal8~0_combout ;
wire \HU|always0~5_combout ;
wire \Mux62~0_combout ;
wire \Mux163~0_combout ;
wire \Mux163~1_combout ;
wire \Mux62~1_combout ;
wire \Mux94~1_combout ;
wire \HU|always0~6_combout ;
wire \HU|ptAScr~4_combout ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \Mux95~0_combout ;
wire \Mux63~0_combout ;
wire \Mux164~0_combout ;
wire \Mux164~1_combout ;
wire \Mux63~1_combout ;
wire \Mux95~1_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux161~0_combout ;
wire \Mux161~1_combout ;
wire \Mux60~0_combout ;
wire \Mux92~0_combout ;
wire \Mux92~1_combout ;
wire \Mux92~2_combout ;
wire \Mux93~0_combout ;
wire \Mux162~0_combout ;
wire \Mux162~1_combout ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \Mux160~0_combout ;
wire \Mux160~1_combout ;
wire \Mux59~0_combout ;
wire \Mux91~0_combout ;
wire \Mux91~1_combout ;
wire \Mux91~2_combout ;
wire \Mux133~0_combout ;
wire \Mux133~1_combout ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \Mux64~0_combout ;
wire \Mux134~0_combout ;
wire \Mux134~1_combout ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \Mux65~0_combout ;
wire \Mux135~0_combout ;
wire \Mux135~1_combout ;
wire \Mux34~0_combout ;
wire \Mux34~1_combout ;
wire \Mux66~0_combout ;
wire \Mux159~0_combout ;
wire \Mux159~1_combout ;
wire \Mux58~0_combout ;
wire \Mux90~2_combout ;
wire \Mux149~0_combout ;
wire \Mux149~1_combout ;
wire \Mux80~2_combout ;
wire \Mux80~3_combout ;
wire \Mux150~0_combout ;
wire \Mux150~1_combout ;
wire \Mux49~0_combout ;
wire \Mux81~2_combout ;
wire \Mux151~0_combout ;
wire \Mux151~1_combout ;
wire \Mux50~0_combout ;
wire \Mux82~2_combout ;
wire \Mux152~0_combout ;
wire \Mux152~1_combout ;
wire \Mux51~0_combout ;
wire \Mux83~2_combout ;
wire \Mux153~0_combout ;
wire \Mux153~1_combout ;
wire \Mux52~0_combout ;
wire \Mux84~2_combout ;
wire \Mux154~0_combout ;
wire \Mux154~1_combout ;
wire \Mux53~0_combout ;
wire \Mux85~2_combout ;
wire \Mux155~0_combout ;
wire \Mux155~1_combout ;
wire \Mux54~0_combout ;
wire \Mux86~2_combout ;
wire \Mux158~0_combout ;
wire \Mux158~1_combout ;
wire \Mux57~0_combout ;
wire \Mux89~3_combout ;
wire \Mux137~0_combout ;
wire \Mux137~1_combout ;
wire \Mux36~0_combout ;
wire \Mux36~1_combout ;
wire \Mux68~0_combout ;
wire \Mux141~0_combout ;
wire \Mux141~1_combout ;
wire \Mux40~0_combout ;
wire \Mux40~1_combout ;
wire \Mux72~0_combout ;
wire \Mux146~0_combout ;
wire \Mux146~1_combout ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \Mux77~0_combout ;
wire \Mux140~0_combout ;
wire \Mux140~1_combout ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \Mux71~0_combout ;
wire \Mux148~0_combout ;
wire \Mux148~1_combout ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \Mux79~0_combout ;
wire \Mux145~0_combout ;
wire \Mux145~1_combout ;
wire \Mux44~0_combout ;
wire \Mux44~1_combout ;
wire \Mux76~0_combout ;
wire \Mux147~0_combout ;
wire \Mux147~1_combout ;
wire \Mux46~0_combout ;
wire \Mux46~1_combout ;
wire \Mux78~0_combout ;
wire \Mux143~0_combout ;
wire \Mux143~1_combout ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \Mux74~0_combout ;
wire \Mux144~0_combout ;
wire \Mux144~1_combout ;
wire \Mux43~0_combout ;
wire \Mux43~1_combout ;
wire \Mux75~0_combout ;
wire \Mux136~0_combout ;
wire \Mux136~1_combout ;
wire \Mux35~0_combout ;
wire \Mux35~1_combout ;
wire \Mux67~0_combout ;
wire \Mux138~0_combout ;
wire \Mux138~1_combout ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \Mux69~0_combout ;
wire \Mux156~0_combout ;
wire \Mux156~1_combout ;
wire \Mux55~0_combout ;
wire \Mux87~2_combout ;
wire \Mux157~0_combout ;
wire \Mux157~1_combout ;
wire \Mux56~0_combout ;
wire \Mux88~2_combout ;
wire \Mux142~0_combout ;
wire \Mux142~1_combout ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \Mux73~0_combout ;
wire \Mux139~0_combout ;
wire \Mux139~1_combout ;
wire \Mux38~0_combout ;
wire \Mux38~1_combout ;
wire \Mux70~0_combout ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Mux93~1_combout ;
wire \Mux93~2_combout ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux4~0_combout ;
wire \Mux4~1_combout ;
wire \ALU|aluif.portOut[1]~15_combout ;
wire \HU|exmem_en~0_combout ;
wire \PR|dmemaddr~0_combout ;
wire \Equal1~0_combout ;
wire \Equal1~1_combout ;
wire \HU|always1~5_combout ;
wire \HU|ifid_en~0_combout ;
wire \PR|dmemren~0_combout ;
wire \PR|dmemwen~0_combout ;
wire \Mux19~2_combout ;
wire \Mux19~3_combout ;
wire \ALU|aluif.portOut[0]~24_combout ;
wire \PR|dmemaddr~1_combout ;
wire \ALU|aluif.portOut[3]~30_combout ;
wire \ALU|aluif.portOut[5]~31_combout ;
wire \ALU|aluif.portOut[2]~33_combout ;
wire \ALU|aluif.portOut[3]~39_combout ;
wire \ALU|aluif.portOut[3]~40_combout ;
wire \PR|dmemaddr~2_combout ;
wire \HU|pc_en~0_combout ;
wire \ALU|aluif.portOut[2]~48_combout ;
wire \PR|dmemaddr~3_combout ;
wire \ALU|aluif.portOut[5]~57_combout ;
wire \ALU|aluif.portOut[5]~58_combout ;
wire \PR|dmemaddr~4_combout ;
wire \ALU|aluif.portOut[4]~65_combout ;
wire \PR|dmemaddr~5_combout ;
wire \ALU|aluif.portOut[7]~72_combout ;
wire \PR|dmemaddr~6_combout ;
wire \ALU|aluif.portOut[6]~79_combout ;
wire \PR|dmemaddr~7_combout ;
wire \ALU|aluif.portOut[9]~90_combout ;
wire \PR|dmemaddr~8_combout ;
wire \ALU|aluif.portOut[8]~96_combout ;
wire \PR|dmemaddr~9_combout ;
wire \ALU|aluif.portOut[11]~102_combout ;
wire \PR|dmemaddr~10_combout ;
wire \ALU|aluif.portOut[10]~108_combout ;
wire \PR|dmemaddr~11_combout ;
wire \ALU|aluif.portOut[13]~114_combout ;
wire \PR|dmemaddr~12_combout ;
wire \ALU|aluif.portOut[12]~120_combout ;
wire \PR|dmemaddr~13_combout ;
wire \ALU|aluif.portOut[15]~126_combout ;
wire \PR|dmemaddr~14_combout ;
wire \ALU|aluif.portOut[14]~132_combout ;
wire \PR|dmemaddr~15_combout ;
wire \ALU|aluif.portOut[23]~140_combout ;
wire \PR|dmemaddr~16_combout ;
wire \ALU|aluif.portOut[22]~147_combout ;
wire \PR|dmemaddr~17_combout ;
wire \ALU|aluif.portOut[21]~153_combout ;
wire \PR|dmemaddr~18_combout ;
wire \ALU|aluif.portOut[29]~166_combout ;
wire \PR|dmemaddr~19_combout ;
wire \ALU|aluif.portOut[28]~180_combout ;
wire \PR|dmemaddr~20_combout ;
wire \ALU|aluif.neg_flag~19_combout ;
wire \PR|dmemaddr~21_combout ;
wire \ALU|aluif.portOut[30]~189_combout ;
wire \PR|dmemaddr~22_combout ;
wire \ALU|aluif.portOut[20]~195_combout ;
wire \PR|dmemaddr~23_combout ;
wire \ALU|aluif.portOut[17]~201_combout ;
wire \PR|dmemaddr~24_combout ;
wire \ALU|aluif.portOut[16]~207_combout ;
wire \PR|dmemaddr~25_combout ;
wire \ALU|aluif.portOut[19]~213_combout ;
wire \PR|dmemaddr~26_combout ;
wire \ALU|aluif.portOut[18]~221_combout ;
wire \PR|dmemaddr~27_combout ;
wire \ALU|aluif.portOut[25]~234_combout ;
wire \PR|dmemaddr~28_combout ;
wire \ALU|aluif.portOut[24]~241_combout ;
wire \PR|dmemaddr~29_combout ;
wire \ALU|aluif.portOut[27]~249_combout ;
wire \PR|dmemaddr~30_combout ;
wire \ALU|aluif.portOut[26]~257_combout ;
wire \PR|dmemaddr~31_combout ;
wire \PR|halt_mem~0_combout ;
wire \PR|dmemstore~0_combout ;
wire \HU|flush_idex~0_combout ;
wire \CU|Equal15~0_combout ;
wire \CU|Equal11~0_combout ;
wire \CU|Equal0~0_combout ;
wire \CU|Equal10~0_combout ;
wire \CU|Equal12~0_combout ;
wire \CU|Equal20~0_combout ;
wire \CU|Equal26~0_combout ;
wire \CU|Equal25~1_combout ;
wire \CU|Equal13~0_combout ;
wire \PR|dataScr_ex~2_combout ;
wire \CU|WideNor0~2_combout ;
wire \CU|Selector0~2_combout ;
wire \PR|ALUOP_ex~0_combout ;
wire \PR|imm_ex~0_combout ;
wire \PR|ALUScr_ex~11_combout ;
wire \PR|shamt_ex~0_combout ;
wire \PR|ALUScr_ex~12_combout ;
wire \PR|Regwen_mem~0_combout ;
wire \PR|regwrite_mem~1_combout ;
wire \PR|regwrite_mem~3_combout ;
wire \PR|regwrite_mem~5_combout ;
wire \PR|regwrite_mem~7_combout ;
wire \PR|regwrite_mem~9_combout ;
wire \PR|rt_ex~0_combout ;
wire \PR|rt_ex~1_combout ;
wire \PR|rt_ex~2_combout ;
wire \PR|rt_ex~3_combout ;
wire \PR|rt_ex~4_combout ;
wire \PR|Regwen_wb~0_combout ;
wire \PR|regwrite_wb~0_combout ;
wire \PR|regwrite_wb~1_combout ;
wire \PR|regwrite_wb~2_combout ;
wire \PR|regwrite_wb~3_combout ;
wire \PR|regwrite_wb~4_combout ;
wire \PR|dmemload_wb~0_combout ;
wire \PR|dmemaddr_wb~0_combout ;
wire \PR|dataScr_wb~0_combout ;
wire \PR|dataScr_wb~1_combout ;
wire \PR|pc_wb~0_combout ;
wire \RF|Mux62~9_combout ;
wire \RF|Mux62~19_combout ;
wire \PR|rdat2_ex~1_combout ;
wire \prif.rs_ex[0]~0_combout ;
wire \PR|prif.rs_ex[1]~0_combout ;
wire \PR|prif.rs_ex[0]~1_combout ;
wire \PR|prif.rs_ex[3]~2_combout ;
wire \PR|prif.rs_ex[2]~3_combout ;
wire \PR|prif.rs_ex[4]~4_combout ;
wire \PR|opcode_mem~0_combout ;
wire \PR|opcode_mem~1_combout ;
wire \PR|opcode_mem~2_combout ;
wire \PR|opcode_mem~3_combout ;
wire \PR|opcode_mem~4_combout ;
wire \PR|opcode_mem~5_combout ;
wire \RF|Mux30~9_combout ;
wire \RF|Mux30~19_combout ;
wire \PR|rdat1_ex~1_combout ;
wire \PR|imm_ex~1_combout ;
wire \PR|shamt_ex~1_combout ;
wire \PR|dmemload_wb~1_combout ;
wire \PR|dmemaddr_wb~1_combout ;
wire \PR|pc_wb~1_combout ;
wire \RF|Mux63~9_combout ;
wire \RF|Mux63~19_combout ;
wire \PR|rdat2_ex~3_combout ;
wire \RF|Mux31~9_combout ;
wire \RF|Mux31~19_combout ;
wire \PR|rdat1_ex~3_combout ;
wire \PR|dmemload_wb~2_combout ;
wire \PR|dmemaddr_wb~2_combout ;
wire \PR|pc_wb~2_combout ;
wire \RF|Mux60~9_combout ;
wire \RF|Mux60~19_combout ;
wire \PR|rdat2_ex~5_combout ;
wire \PR|imm_ex~2_combout ;
wire \PR|shamt_ex~2_combout ;
wire \PR|imm_ex~3_combout ;
wire \PR|shamt_ex~3_combout ;
wire \PR|dmemload_wb~3_combout ;
wire \PR|dmemaddr_wb~3_combout ;
wire \PR|pc_wb~3_combout ;
wire \RF|Mux61~9_combout ;
wire \RF|Mux61~19_combout ;
wire \PR|rdat2_ex~7_combout ;
wire \PR|dmemload_wb~4_combout ;
wire \PR|dmemaddr_wb~4_combout ;
wire \PR|pc_wb~4_combout ;
wire \RF|Mux59~9_combout ;
wire \RF|Mux59~19_combout ;
wire \PR|rdat2_ex~9_combout ;
wire \PR|imm_ex~4_combout ;
wire \PR|shamt_ex~4_combout ;
wire \PR|instr_ex~0_combout ;
wire \PR|dmemload_wb~5_combout ;
wire \PR|imm_wb~0_combout ;
wire \PR|dmemaddr_wb~5_combout ;
wire \PR|pc_wb~5_combout ;
wire \RF|Mux32~9_combout ;
wire \RF|Mux32~19_combout ;
wire \PR|rdat2_ex~11_combout ;
wire \PR|imm_mem~0_combout ;
wire \PR|imm_wb~1_combout ;
wire \PR|dmemload_wb~6_combout ;
wire \PR|dmemaddr_wb~6_combout ;
wire \PR|pc_wb~6_combout ;
wire \RF|Mux33~9_combout ;
wire \RF|Mux33~19_combout ;
wire \PR|rdat2_ex~13_combout ;
wire \PR|imm_mem~1_combout ;
wire \PR|dmemload_wb~7_combout ;
wire \PR|imm_wb~2_combout ;
wire \PR|dmemaddr_wb~7_combout ;
wire \PR|pc_wb~7_combout ;
wire \RF|Mux34~9_combout ;
wire \RF|Mux34~19_combout ;
wire \PR|rdat2_ex~15_combout ;
wire \PR|imm_mem~2_combout ;
wire \PR|imm_ex~5_combout ;
wire \PR|dmemload_wb~8_combout ;
wire \PR|dmemaddr_wb~8_combout ;
wire \PR|pc_wb~8_combout ;
wire \RF|Mux58~9_combout ;
wire \RF|Mux58~19_combout ;
wire \PR|rdat2_ex~17_combout ;
wire \PR|imm_ex~6_combout ;
wire \PR|dmemload_wb~9_combout ;
wire \PR|dmemaddr_wb~9_combout ;
wire \PR|pc_wb~9_combout ;
wire \RF|Mux48~9_combout ;
wire \RF|Mux48~19_combout ;
wire \PR|rdat2_ex~19_combout ;
wire \PR|imm_ex~7_combout ;
wire \PR|dmemload_wb~10_combout ;
wire \PR|dmemaddr_wb~10_combout ;
wire \PR|pc_wb~10_combout ;
wire \RF|Mux49~9_combout ;
wire \RF|Mux49~19_combout ;
wire \PR|rdat2_ex~21_combout ;
wire \PR|imm_ex~8_combout ;
wire \PR|dmemload_wb~11_combout ;
wire \PR|dmemaddr_wb~11_combout ;
wire \PR|pc_wb~11_combout ;
wire \RF|Mux50~9_combout ;
wire \RF|Mux50~19_combout ;
wire \PR|rdat2_ex~23_combout ;
wire \PR|imm_ex~9_combout ;
wire \PR|dmemload_wb~12_combout ;
wire \PR|dmemaddr_wb~12_combout ;
wire \PR|pc_wb~12_combout ;
wire \RF|Mux51~9_combout ;
wire \RF|Mux51~19_combout ;
wire \PR|rdat2_ex~25_combout ;
wire \PR|imm_ex~10_combout ;
wire \PR|dmemload_wb~13_combout ;
wire \PR|dmemaddr_wb~13_combout ;
wire \PR|pc_wb~13_combout ;
wire \RF|Mux52~9_combout ;
wire \RF|Mux52~19_combout ;
wire \PR|rdat2_ex~27_combout ;
wire \PR|imm_ex~11_combout ;
wire \PR|dmemload_wb~14_combout ;
wire \PR|dmemaddr_wb~14_combout ;
wire \PR|pc_wb~14_combout ;
wire \RF|Mux53~9_combout ;
wire \RF|Mux53~19_combout ;
wire \PR|rdat2_ex~29_combout ;
wire \PR|imm_ex~12_combout ;
wire \PR|dmemload_wb~15_combout ;
wire \PR|dmemaddr_wb~15_combout ;
wire \PR|pc_wb~15_combout ;
wire \RF|Mux54~9_combout ;
wire \RF|Mux54~19_combout ;
wire \PR|rdat2_ex~31_combout ;
wire \PR|imm_ex~13_combout ;
wire \PR|dmemload_wb~16_combout ;
wire \PR|dmemaddr_wb~16_combout ;
wire \PR|pc_wb~16_combout ;
wire \RF|Mux57~9_combout ;
wire \RF|Mux57~19_combout ;
wire \PR|rdat2_ex~33_combout ;
wire \PR|dmemload_wb~17_combout ;
wire \PR|imm_wb~3_combout ;
wire \PR|dmemaddr_wb~17_combout ;
wire \PR|pc_wb~17_combout ;
wire \RF|Mux36~9_combout ;
wire \RF|Mux36~19_combout ;
wire \PR|rdat2_ex~35_combout ;
wire \PR|imm_mem~3_combout ;
wire \PR|dmemload_wb~18_combout ;
wire \PR|imm_wb~4_combout ;
wire \PR|dmemaddr_wb~18_combout ;
wire \PR|pc_wb~18_combout ;
wire \RF|Mux40~9_combout ;
wire \RF|Mux40~19_combout ;
wire \PR|rdat2_ex~37_combout ;
wire \PR|imm_mem~4_combout ;
wire \PR|imm_wb~5_combout ;
wire \PR|dmemload_wb~19_combout ;
wire \PR|dmemaddr_wb~19_combout ;
wire \PR|pc_wb~19_combout ;
wire \RF|Mux45~9_combout ;
wire \RF|Mux45~19_combout ;
wire \PR|rdat2_ex~39_combout ;
wire \PR|imm_mem~5_combout ;
wire \PR|imm_wb~6_combout ;
wire \PR|dmemload_wb~20_combout ;
wire \PR|dmemaddr_wb~20_combout ;
wire \PR|pc_wb~20_combout ;
wire \RF|Mux39~9_combout ;
wire \RF|Mux39~19_combout ;
wire \PR|rdat2_ex~41_combout ;
wire \PR|imm_mem~6_combout ;
wire \PR|imm_wb~7_combout ;
wire \PR|dmemload_wb~21_combout ;
wire \PR|dmemaddr_wb~21_combout ;
wire \PR|pc_wb~21_combout ;
wire \RF|Mux47~9_combout ;
wire \RF|Mux47~19_combout ;
wire \PR|rdat2_ex~43_combout ;
wire \PR|imm_mem~7_combout ;
wire \PR|dmemload_wb~22_combout ;
wire \PR|imm_wb~8_combout ;
wire \PR|dmemaddr_wb~22_combout ;
wire \PR|pc_wb~22_combout ;
wire \RF|Mux44~9_combout ;
wire \RF|Mux44~19_combout ;
wire \PR|rdat2_ex~45_combout ;
wire \PR|imm_mem~8_combout ;
wire \PR|dmemload_wb~23_combout ;
wire \PR|imm_wb~9_combout ;
wire \PR|dmemaddr_wb~23_combout ;
wire \PR|pc_wb~23_combout ;
wire \RF|Mux46~9_combout ;
wire \RF|Mux46~19_combout ;
wire \PR|rdat2_ex~47_combout ;
wire \PR|imm_mem~9_combout ;
wire \PR|dmemload_wb~24_combout ;
wire \PR|imm_wb~10_combout ;
wire \PR|dmemaddr_wb~24_combout ;
wire \PR|pc_wb~24_combout ;
wire \RF|Mux42~9_combout ;
wire \RF|Mux42~19_combout ;
wire \PR|rdat2_ex~49_combout ;
wire \PR|imm_mem~10_combout ;
wire \PR|imm_wb~11_combout ;
wire \PR|dmemload_wb~25_combout ;
wire \PR|dmemaddr_wb~25_combout ;
wire \PR|pc_wb~25_combout ;
wire \RF|Mux43~9_combout ;
wire \RF|Mux43~19_combout ;
wire \PR|rdat2_ex~51_combout ;
wire \PR|imm_mem~11_combout ;
wire \PR|imm_wb~12_combout ;
wire \PR|dmemload_wb~26_combout ;
wire \PR|dmemaddr_wb~26_combout ;
wire \PR|pc_wb~26_combout ;
wire \RF|Mux35~9_combout ;
wire \RF|Mux35~19_combout ;
wire \PR|rdat2_ex~53_combout ;
wire \PR|imm_mem~12_combout ;
wire \PR|imm_wb~13_combout ;
wire \PR|dmemload_wb~27_combout ;
wire \PR|dmemaddr_wb~27_combout ;
wire \PR|pc_wb~27_combout ;
wire \RF|Mux37~9_combout ;
wire \RF|Mux37~19_combout ;
wire \PR|rdat2_ex~55_combout ;
wire \PR|imm_mem~13_combout ;
wire \PR|imm_ex~14_combout ;
wire \PR|dmemload_wb~28_combout ;
wire \PR|dmemaddr_wb~28_combout ;
wire \PR|pc_wb~28_combout ;
wire \RF|Mux55~9_combout ;
wire \RF|Mux55~19_combout ;
wire \PR|rdat2_ex~57_combout ;
wire \PR|imm_ex~15_combout ;
wire \PR|dmemload_wb~29_combout ;
wire \PR|dmemaddr_wb~29_combout ;
wire \PR|pc_wb~29_combout ;
wire \RF|Mux56~9_combout ;
wire \RF|Mux56~19_combout ;
wire \PR|rdat2_ex~59_combout ;
wire \PR|imm_wb~14_combout ;
wire \PR|dmemload_wb~30_combout ;
wire \PR|dmemaddr_wb~30_combout ;
wire \PR|pc_wb~30_combout ;
wire \RF|Mux41~9_combout ;
wire \RF|Mux41~19_combout ;
wire \PR|rdat2_ex~61_combout ;
wire \PR|imm_mem~14_combout ;
wire \PR|dmemload_wb~31_combout ;
wire \PR|imm_wb~15_combout ;
wire \PR|dmemaddr_wb~31_combout ;
wire \PR|pc_wb~31_combout ;
wire \RF|Mux38~9_combout ;
wire \RF|Mux38~19_combout ;
wire \PR|rdat2_ex~63_combout ;
wire \PR|imm_mem~15_combout ;
wire \CU|Equal4~0_combout ;
wire \PR|ALUOP_ex~2_combout ;
wire \CU|Selector2~4_combout ;
wire \CU|Selector2~5_combout ;
wire \PR|ALUOP_ex~3_combout ;
wire \RF|Mux29~9_combout ;
wire \RF|Mux29~19_combout ;
wire \PR|rdat1_ex~5_combout ;
wire \RF|Mux27~9_combout ;
wire \RF|Mux27~19_combout ;
wire \PR|rdat1_ex~7_combout ;
wire \RF|Mux28~9_combout ;
wire \RF|Mux28~19_combout ;
wire \PR|rdat1_ex~9_combout ;
wire \RF|Mux23~9_combout ;
wire \RF|Mux23~19_combout ;
wire \PR|rdat1_ex~11_combout ;
wire \RF|Mux24~9_combout ;
wire \RF|Mux24~19_combout ;
wire \PR|rdat1_ex~13_combout ;
wire \RF|Mux25~9_combout ;
wire \RF|Mux25~19_combout ;
wire \PR|rdat1_ex~15_combout ;
wire \RF|Mux26~9_combout ;
wire \RF|Mux26~19_combout ;
wire \PR|rdat1_ex~17_combout ;
wire \RF|Mux15~9_combout ;
wire \RF|Mux15~19_combout ;
wire \PR|rdat1_ex~19_combout ;
wire \RF|Mux16~9_combout ;
wire \RF|Mux16~19_combout ;
wire \PR|rdat1_ex~21_combout ;
wire \RF|Mux17~9_combout ;
wire \RF|Mux17~19_combout ;
wire \PR|rdat1_ex~23_combout ;
wire \RF|Mux18~9_combout ;
wire \RF|Mux18~19_combout ;
wire \PR|rdat1_ex~25_combout ;
wire \RF|Mux20~9_combout ;
wire \RF|Mux20~19_combout ;
wire \PR|rdat1_ex~27_combout ;
wire \RF|Mux19~9_combout ;
wire \RF|Mux19~19_combout ;
wire \PR|rdat1_ex~29_combout ;
wire \RF|Mux21~9_combout ;
wire \RF|Mux21~19_combout ;
wire \PR|rdat1_ex~31_combout ;
wire \RF|Mux22~9_combout ;
wire \RF|Mux22~19_combout ;
wire \PR|rdat1_ex~33_combout ;
wire \RF|Mux13~9_combout ;
wire \RF|Mux13~19_combout ;
wire \PR|rdat1_ex~35_combout ;
wire \RF|Mux14~9_combout ;
wire \RF|Mux14~19_combout ;
wire \PR|rdat1_ex~37_combout ;
wire \RF|Mux11~9_combout ;
wire \RF|Mux11~19_combout ;
wire \PR|rdat1_ex~39_combout ;
wire \RF|Mux12~9_combout ;
wire \RF|Mux12~19_combout ;
wire \PR|rdat1_ex~41_combout ;
wire \RF|Mux9~9_combout ;
wire \RF|Mux9~19_combout ;
wire \PR|rdat1_ex~43_combout ;
wire \RF|Mux10~9_combout ;
wire \RF|Mux10~19_combout ;
wire \PR|rdat1_ex~45_combout ;
wire \RF|Mux7~9_combout ;
wire \RF|Mux7~19_combout ;
wire \PR|rdat1_ex~47_combout ;
wire \RF|Mux8~9_combout ;
wire \RF|Mux8~19_combout ;
wire \PR|rdat1_ex~49_combout ;
wire \RF|Mux0~9_combout ;
wire \RF|Mux0~19_combout ;
wire \PR|rdat1_ex~51_combout ;
wire \RF|Mux1~9_combout ;
wire \RF|Mux1~19_combout ;
wire \PR|rdat1_ex~53_combout ;
wire \RF|Mux2~9_combout ;
wire \RF|Mux2~19_combout ;
wire \PR|rdat1_ex~55_combout ;
wire \RF|Mux5~9_combout ;
wire \RF|Mux5~19_combout ;
wire \PR|rdat1_ex~57_combout ;
wire \RF|Mux6~9_combout ;
wire \RF|Mux6~19_combout ;
wire \PR|rdat1_ex~59_combout ;
wire \RF|Mux3~9_combout ;
wire \RF|Mux3~19_combout ;
wire \PR|rdat1_ex~61_combout ;
wire \RF|Mux4~9_combout ;
wire \RF|Mux4~19_combout ;
wire \PR|rdat1_ex~63_combout ;
wire \PR|ALUScr_ex~13_combout ;
wire \CU|Selector3~5_combout ;
wire \PR|ALUOP_ex~4_combout ;
wire \ALU|aluif.portOut[5]~258_combout ;
wire \PR|instr_mem~0_combout ;
wire \PR|instr_mem~1_combout ;
wire \PR|instr_mem~2_combout ;
wire \PR|instr_mem~3_combout ;
wire \PR|instr_mem~4_combout ;
wire \PR|instr_mem~5_combout ;
wire \PR|rdat1_mem~0_combout ;
wire \PR|PCScr_mem~0_combout ;
wire \PR|pc_bran_mem~0_combout ;
wire \PR|PCScr_mem~1_combout ;
wire \PR|opcode_ex~0_combout ;
wire \PR|opcode_ex~1_combout ;
wire \PR|opcode_ex~2_combout ;
wire \PR|opcode_ex~3_combout ;
wire \PR|opcode_ex~4_combout ;
wire \CU|Equal13~1_combout ;
wire \PR|memren_ex~0_combout ;
wire \PR|memwen_ex~0_combout ;
wire \PR|rdat1_mem~1_combout ;
wire \PR|pc_bran_mem~1_combout ;
wire \PR|rdat1_mem~2_combout ;
wire \PR|pc_bran_mem~2_combout ;
wire \PR|rdat1_mem~3_combout ;
wire \PR|pc_bran_mem~3_combout ;
wire \PR|rdat1_mem~4_combout ;
wire \PR|pc_bran_mem~4_combout ;
wire \PR|rdat1_mem~5_combout ;
wire \PR|pc_bran_mem~5_combout ;
wire \PR|rdat1_mem~6_combout ;
wire \PR|pc_bran_mem~6_combout ;
wire \PR|rdat1_mem~7_combout ;
wire \PR|pc_bran_mem~7_combout ;
wire \PR|rdat1_mem~8_combout ;
wire \PR|pc_bran_mem~8_combout ;
wire \PR|instr_mem~6_combout ;
wire \PR|rdat1_mem~9_combout ;
wire \PR|pc_bran_mem~9_combout ;
wire \PR|instr_mem~7_combout ;
wire \PR|rdat1_mem~10_combout ;
wire \PR|pc_bran_mem~10_combout ;
wire \PR|instr_mem~8_combout ;
wire \PR|rdat1_mem~11_combout ;
wire \PR|pc_bran_mem~11_combout ;
wire \PR|instr_mem~9_combout ;
wire \PR|rdat1_mem~12_combout ;
wire \PR|pc_bran_mem~12_combout ;
wire \PR|instr_mem~10_combout ;
wire \PR|rdat1_mem~13_combout ;
wire \PR|pc_bran_mem~13_combout ;
wire \PR|instr_mem~11_combout ;
wire \PR|rdat1_mem~14_combout ;
wire \PR|pc_bran_mem~14_combout ;
wire \PR|instr_mem~12_combout ;
wire \PR|rdat1_mem~15_combout ;
wire \PR|pc_bran_mem~15_combout ;
wire \PR|instr_mem~13_combout ;
wire \PR|rdat1_mem~16_combout ;
wire \PR|pc_bran_mem~16_combout ;
wire \PR|instr_mem~14_combout ;
wire \PR|rdat1_mem~17_combout ;
wire \PR|pc_bran_mem~17_combout ;
wire \PR|instr_mem~15_combout ;
wire \PR|rdat1_mem~18_combout ;
wire \PR|pc_bran_mem~18_combout ;
wire \PR|instr_mem~16_combout ;
wire \PR|rdat1_mem~19_combout ;
wire \PR|pc_bran_mem~19_combout ;
wire \prif.pc_mem[15]~0_combout ;
wire \PR|prif.pc_mem[29]~0_combout ;
wire \PR|rdat1_mem~20_combout ;
wire \PR|pc_bran_mem~20_combout ;
wire \PR|prif.pc_mem[28]~1_combout ;
wire \PR|rdat1_mem~21_combout ;
wire \PR|pc_bran_mem~21_combout ;
wire \PR|prif.pc_mem[31]~2_combout ;
wire \PR|rdat1_mem~22_combout ;
wire \PR|pc_bran_mem~22_combout ;
wire \PR|prif.pc_mem[30]~3_combout ;
wire \PR|rdat1_mem~23_combout ;
wire \PR|pc_bran_mem~23_combout ;
wire \PR|instr_mem~17_combout ;
wire \PR|rdat1_mem~24_combout ;
wire \PR|pc_bran_mem~24_combout ;
wire \PR|instr_mem~18_combout ;
wire \PR|rdat1_mem~25_combout ;
wire \PR|pc_bran_mem~25_combout ;
wire \PR|instr_mem~19_combout ;
wire \PR|rdat1_mem~26_combout ;
wire \PR|pc_bran_mem~26_combout ;
wire \PR|instr_mem~20_combout ;
wire \PR|rdat1_mem~27_combout ;
wire \PR|pc_bran_mem~27_combout ;
wire \PR|instr_mem~21_combout ;
wire \PR|rdat1_mem~28_combout ;
wire \PR|pc_bran_mem~28_combout ;
wire \PR|instr_mem~22_combout ;
wire \PR|rdat1_mem~29_combout ;
wire \PR|pc_bran_mem~29_combout ;
wire \PR|instr_mem~23_combout ;
wire \PR|rdat1_mem~30_combout ;
wire \PR|pc_bran_mem~30_combout ;
wire \PR|instr_mem~24_combout ;
wire \PR|rdat1_mem~31_combout ;
wire \PR|pc_bran_mem~31_combout ;
wire \PR|instr_mem~25_combout ;
wire \PR|dmemstore~1_combout ;
wire \PR|dmemstore~2_combout ;
wire \Mux60~1_combout ;
wire \PR|dmemstore~3_combout ;
wire \Mux59~1_combout ;
wire \PR|dmemstore~4_combout ;
wire \Mux58~1_combout ;
wire \PR|dmemstore~5_combout ;
wire \Mux57~1_combout ;
wire \PR|dmemstore~6_combout ;
wire \Mux56~1_combout ;
wire \PR|dmemstore~7_combout ;
wire \Mux55~1_combout ;
wire \PR|dmemstore~8_combout ;
wire \Mux54~1_combout ;
wire \PR|dmemstore~9_combout ;
wire \Mux53~1_combout ;
wire \PR|dmemstore~10_combout ;
wire \Mux52~1_combout ;
wire \PR|dmemstore~11_combout ;
wire \Mux51~1_combout ;
wire \PR|dmemstore~12_combout ;
wire \Mux50~1_combout ;
wire \PR|dmemstore~13_combout ;
wire \Mux49~1_combout ;
wire \PR|dmemstore~14_combout ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \PR|dmemstore~15_combout ;
wire \PR|dmemstore~16_combout ;
wire \PR|dmemstore~17_combout ;
wire \PR|dmemstore~18_combout ;
wire \PR|dmemstore~19_combout ;
wire \PR|dmemstore~20_combout ;
wire \PR|dmemstore~21_combout ;
wire \PR|dmemstore~22_combout ;
wire \PR|dmemstore~23_combout ;
wire \PR|dmemstore~24_combout ;
wire \PR|dmemstore~25_combout ;
wire \PR|dmemstore~26_combout ;
wire \PR|dmemstore~27_combout ;
wire \PR|dmemstore~28_combout ;
wire \PR|dmemstore~29_combout ;
wire \PR|dmemstore~30_combout ;
wire \PR|dmemstore~31_combout ;
wire \PR|halt_ex~0_combout ;
wire \prif.halt_wb~q ;
wire \HU|ifid_en~1_combout ;
wire \PR|imemload_id~0_combout ;
wire \PR|imemload_id~1_combout ;
wire \PR|imemload_id~2_combout ;
wire \PR|imemload_id~3_combout ;
wire \PR|imemload_id~4_combout ;
wire \PR|imemload_id~5_combout ;
wire \PR|imemload_id~6_combout ;
wire \PR|imemload_id~7_combout ;
wire \PR|imemload_id~8_combout ;
wire \PR|imemload_id~9_combout ;
wire \PR|imemload_id~10_combout ;
wire \PR|imemload_id~11_combout ;
wire \PR|imemload_id~12_combout ;
wire \PR|Regwen_ex~0_combout ;
wire \PR|rd_ex~0_combout ;
wire \PR|RegDest_ex~0_combout ;
wire \PR|RegDest_ex~1_combout ;
wire \PR|rd_ex~1_combout ;
wire \PR|rd_ex~2_combout ;
wire \PR|rd_ex~3_combout ;
wire \PR|rd_ex~4_combout ;
wire \PR|imemload_id~13_combout ;
wire \PR|imemload_id~14_combout ;
wire \PR|imemload_id~15_combout ;
wire \PR|imemload_id~16_combout ;
wire \PR|imemload_id~17_combout ;
wire \PR|dataScr_mem~0_combout ;
wire \PR|dataScr_mem~1_combout ;
wire \PR|prif.pc_mem[1]~4_combout ;
wire \PR|imemload_id~18_combout ;
wire \PR|imemload_id~19_combout ;
wire \PR|imemload_id~20_combout ;
wire \PR|imemload_id~21_combout ;
wire \PR|imemload_id~22_combout ;
wire \PR|opcode_ex~5_combout ;
wire \PR|imemload_id~23_combout ;
wire \PR|prif.pc_mem[0]~5_combout ;
wire \PR|prif.pc_mem[3]~6_combout ;
wire \PR|imemload_id~24_combout ;
wire \PR|imemload_id~25_combout ;
wire \PR|prif.pc_mem[2]~7_combout ;
wire \PR|prif.pc_mem[4]~8_combout ;
wire \PR|imemload_id~26_combout ;
wire \PR|imemload_id~27_combout ;
wire \PR|prif.pc_mem[5]~9_combout ;
wire \PR|prif.pc_mem[15]~10_combout ;
wire \PR|imemload_id~28_combout ;
wire \PR|prif.pc_mem[14]~11_combout ;
wire \PR|imemload_id~29_combout ;
wire \PR|prif.pc_mem[13]~12_combout ;
wire \PR|imemload_id~30_combout ;
wire \PR|prif.pc_mem[12]~13_combout ;
wire \PR|imemload_id~31_combout ;
wire \PR|prif.pc_mem[11]~14_combout ;
wire \PR|prif.pc_mem[10]~15_combout ;
wire \PR|prif.pc_mem[9]~16_combout ;
wire \PR|prif.pc_mem[6]~17_combout ;
wire \PR|prif.pc_mem[27]~18_combout ;
wire \PR|prif.pc_mem[23]~19_combout ;
wire \PR|prif.pc_mem[18]~20_combout ;
wire \PR|prif.pc_mem[24]~21_combout ;
wire \PR|prif.pc_mem[16]~22_combout ;
wire \PR|prif.pc_mem[19]~23_combout ;
wire \PR|prif.pc_mem[17]~24_combout ;
wire \PR|prif.pc_mem[21]~25_combout ;
wire \PR|prif.pc_mem[20]~26_combout ;
wire \PR|prif.pc_mem[26]~27_combout ;
wire \PR|prif.pc_mem[8]~28_combout ;
wire \PR|prif.pc_mem[7]~29_combout ;
wire \PR|prif.pc_mem[22]~30_combout ;
wire \PR|prif.pc_mem[25]~31_combout ;
wire \PR|instr_ex~1_combout ;
wire \PR|instr_ex~2_combout ;
wire \PR|instr_ex~3_combout ;
wire \PR|instr_ex~4_combout ;
wire \PR|instr_ex~5_combout ;
wire \PR|instr_ex~6_combout ;
wire \PR|PCScr_ex~3_combout ;
wire \PR|pc_ex~0_combout ;
wire \PR|PCScr_ex~4_combout ;
wire \PR|pc_ex~1_combout ;
wire \PR|pc_ex~2_combout ;
wire \PR|pc_ex~3_combout ;
wire \PR|pc_ex~4_combout ;
wire \PR|pc_ex~5_combout ;
wire \PR|pc_ex~6_combout ;
wire \PR|pc_ex~7_combout ;
wire \PR|pc_ex~8_combout ;
wire \PR|pc_ex~9_combout ;
wire \PR|instr_ex~7_combout ;
wire \PR|instr_ex~8_combout ;
wire \PR|pc_ex~10_combout ;
wire \PR|pc_ex~11_combout ;
wire \PR|instr_ex~9_combout ;
wire \PR|instr_ex~10_combout ;
wire \PR|pc_ex~12_combout ;
wire \PR|pc_ex~13_combout ;
wire \PR|instr_ex~11_combout ;
wire \PR|instr_ex~12_combout ;
wire \PR|pc_ex~14_combout ;
wire \PR|pc_ex~15_combout ;
wire \PR|instr_ex~13_combout ;
wire \PR|instr_ex~14_combout ;
wire \PR|pc_ex~16_combout ;
wire \PR|pc_ex~17_combout ;
wire \PR|pc_ex~18_combout ;
wire \PR|pc_ex~19_combout ;
wire \PR|pc_ex~20_combout ;
wire \PR|pc_ex~21_combout ;
wire \PR|pc_ex~22_combout ;
wire \PR|pc_ex~23_combout ;
wire \PR|instr_ex~15_combout ;
wire \PR|instr_ex~16_combout ;
wire \PR|instr_ex~17_combout ;
wire \PR|pc_ex~24_combout ;
wire \PR|pc_ex~25_combout ;
wire \PR|pc_ex~26_combout ;
wire \PR|pc_ex~27_combout ;
wire \PR|pc_ex~28_combout ;
wire \PR|pc_ex~29_combout ;
wire \PR|pc_ex~30_combout ;
wire \PR|pc_ex~31_combout ;
wire \PR|instr_ex~18_combout ;
wire \PR|instr_ex~19_combout ;
wire \PR|instr_ex~20_combout ;
wire \PR|instr_ex~21_combout ;
wire \PR|instr_ex~22_combout ;
wire \PR|instr_ex~23_combout ;
wire \PR|instr_ex~24_combout ;
wire \PR|instr_ex~25_combout ;
wire \PR|halt_wb~0_combout ;
wire \PR|dataScr_ex~3_combout ;
wire \PR|pc_id~0_combout ;
wire \PR|pc_id~1_combout ;
wire \PR|pc_id~2_combout ;
wire \PR|pc_id~3_combout ;
wire \PR|pc_id~4_combout ;
wire \PR|pc_id~5_combout ;
wire \PR|pc_id~6_combout ;
wire \PR|pc_id~7_combout ;
wire \PR|pc_id~8_combout ;
wire \PR|pc_id~9_combout ;
wire \PR|pc_id~10_combout ;
wire \PR|pc_id~11_combout ;
wire \PR|pc_id~12_combout ;
wire \PR|pc_id~13_combout ;
wire \PR|pc_id~14_combout ;
wire \PR|pc_id~15_combout ;
wire \PR|pc_id~16_combout ;
wire \PR|pc_id~17_combout ;
wire \PR|pc_id~18_combout ;
wire \PR|pc_id~19_combout ;
wire \PR|pc_id~20_combout ;
wire \PR|pc_id~21_combout ;
wire \PR|pc_id~22_combout ;
wire \PR|pc_id~23_combout ;
wire \PR|pc_id~24_combout ;
wire \PR|pc_id~25_combout ;
wire \PR|pc_id~26_combout ;
wire \PR|pc_id~27_combout ;
wire \PR|pc_id~28_combout ;
wire \PR|pc_id~29_combout ;
wire \PR|pc_id~30_combout ;
wire \PR|pc_id~31_combout ;
wire \Mux90~3_combout ;
wire \Mux80~4_combout ;
wire \Mux81~3_combout ;
wire \Mux82~3_combout ;
wire \Mux83~3_combout ;
wire \Mux84~3_combout ;
wire \Mux85~3_combout ;
wire \Mux86~3_combout ;
wire \Mux89~4_combout ;
wire \Mux87~3_combout ;
wire \Mux88~3_combout ;
wire \PR|dataScr_ex~4_combout ;
wire \PR|ALUScr_ex~15_combout ;
wire \PR|zero_flag_mem~13_combout ;
wire \prif.ALUScr_ex[0]~feeder_combout ;
wire \prif.rdat1_mem[21]~0_combout ;
wire \Mux131~0_combout ;
wire \prif.zero_flag_mem~q ;
wire \pc[0]~0_combout ;
wire \pc[1]~1_combout ;
wire \Mux132~0_combout ;
wire \pc[23]~2_combout ;
wire \Add3~1 ;
wire \Add3~2_combout ;
wire \Mux129~0_combout ;
wire \Mux129~1_combout ;
wire \Mux130~0_combout ;
wire \Add3~0_combout ;
wire \Mux130~1_combout ;
wire \Add3~3 ;
wire \Add3~5 ;
wire \Add3~6_combout ;
wire \Mux127~0_combout ;
wire \Mux127~1_combout ;
wire \Mux128~0_combout ;
wire \Add3~4_combout ;
wire \Mux128~1_combout ;
wire \Add3~7 ;
wire \Add3~9 ;
wire \Add3~10_combout ;
wire \Mux125~0_combout ;
wire \Mux125~1_combout ;
wire \Mux126~0_combout ;
wire \Add3~8_combout ;
wire \Mux126~1_combout ;
wire \Mux123~0_combout ;
wire \Mux123~1_combout ;
wire \Add3~11 ;
wire \Add3~12_combout ;
wire \Mux124~0_combout ;
wire \Mux124~1_combout ;
wire \Add3~13 ;
wire \Add3~15 ;
wire \Add3~17 ;
wire \Add3~18_combout ;
wire \Mux121~0_combout ;
wire \Mux121~1_combout ;
wire \Mux122~0_combout ;
wire \Add3~16_combout ;
wire \Mux122~1_combout ;
wire \Add3~19 ;
wire \Add3~21 ;
wire \Add3~22_combout ;
wire \Mux119~0_combout ;
wire \Mux119~1_combout ;
wire \Add3~20_combout ;
wire \Mux120~0_combout ;
wire \Mux120~1_combout ;
wire \Add3~23 ;
wire \Add3~25 ;
wire \Add3~26_combout ;
wire \Mux117~0_combout ;
wire \Mux117~1_combout ;
wire \Add3~24_combout ;
wire \Mux118~0_combout ;
wire \Mux118~1_combout ;
wire \Add3~27 ;
wire \Add3~29 ;
wire \Add3~31 ;
wire \Add3~33 ;
wire \Add3~35 ;
wire \Add3~37 ;
wire \Add3~39 ;
wire \Add3~41 ;
wire \Add3~42_combout ;
wire \Mux109~0_combout ;
wire \Mux109~1_combout ;
wire \Mux110~0_combout ;
wire \Add3~40_combout ;
wire \Mux110~1_combout ;
wire \Add3~38_combout ;
wire \Mux111~0_combout ;
wire \Mux111~1_combout ;
wire \Mux103~0_combout ;
wire \Add3~43 ;
wire \Add3~45 ;
wire \Add3~47 ;
wire \Add3~49 ;
wire \Add3~51 ;
wire \Add3~53 ;
wire \Add3~54_combout ;
wire \Mux103~1_combout ;
wire \Add3~52_combout ;
wire \Mux104~0_combout ;
wire \Mux104~1_combout ;
wire \Add3~55 ;
wire \Add3~57 ;
wire \Add3~58_combout ;
wire \Mux101~0_combout ;
wire \Mux101~1_combout ;
wire \Add3~56_combout ;
wire \Mux102~0_combout ;
wire \Mux102~1_combout ;
wire \Add3~36_combout ;
wire \Mux112~0_combout ;
wire \Mux112~1_combout ;
wire \Mux115~0_combout ;
wire \Mux115~1_combout ;
wire \Add3~28_combout ;
wire \Mux116~0_combout ;
wire \Mux116~1_combout ;
wire \Mux113~0_combout ;
wire \Mux113~1_combout ;
wire \Mux114~0_combout ;
wire \Add3~32_combout ;
wire \Mux114~1_combout ;
wire \Mux107~0_combout ;
wire \Mux107~1_combout ;
wire \Add3~44_combout ;
wire \Mux108~0_combout ;
wire \Mux108~1_combout ;
wire \Add3~50_combout ;
wire \Mux105~0_combout ;
wire \Mux105~1_combout ;
wire \Mux106~0_combout ;
wire \Add3~48_combout ;
wire \Mux106~1_combout ;
wire \dpif.halt~_Duplicate_1_q ;
wire \prif.halt_mem~q ;
wire \dpif.halt~0_combout ;
wire [4:0] \prif.shamt_ex ;
wire [4:0] \prif.rt_ex ;
wire [4:0] \prif.rs_ex ;
wire [4:0] \prif.regwrite_wb ;
wire [4:0] \prif.regwrite_mem ;
wire [31:0] \prif.rdat2_ex ;
wire [31:0] \prif.rdat1_mem ;
wire [31:0] \prif.rdat1_ex ;
wire [4:0] \prif.rd_ex ;
wire [31:0] \prif.pc_wb ;
wire [31:0] \prif.pc_mem ;
wire [31:0] \prif.pc_id ;
wire [31:0] \prif.pc_ex ;
wire [31:0] \prif.pc_bran_mem ;
wire [5:0] \prif.opcode_mem ;
wire [5:0] \prif.opcode_ex ;
wire [31:0] \prif.instr_mem ;
wire [31:0] \prif.instr_ex ;
wire [15:0] \prif.imm_wb ;
wire [15:0] \prif.imm_mem ;
wire [15:0] \prif.imm_ex ;
wire [31:0] \prif.imemload_id ;
wire [31:0] \prif.dmemload_wb ;
wire [31:0] \prif.dmemaddr_wb ;
wire [1:0] \prif.dataScr_wb ;
wire [1:0] \prif.dataScr_mem ;
wire [1:0] \prif.dataScr_ex ;
wire [1:0] \prif.RegDest_ex ;
wire [1:0] \prif.PCScr_mem ;
wire [1:0] \prif.PCScr_ex ;
wire [1:0] \prif.ALUScr_ex ;
wire [3:0] \prif.ALUOP_ex ;


hazard_unit HU(
	.prifRegwen_mem(\prif.Regwen_mem~q ),
	.prifregwrite_mem_4(\prif.regwrite_mem [4]),
	.prifregwrite_mem_0(\prif.regwrite_mem [0]),
	.prifregwrite_mem_1(\prif.regwrite_mem [1]),
	.prifregwrite_mem_2(\prif.regwrite_mem [2]),
	.prifregwrite_mem_3(\prif.regwrite_mem [3]),
	.prifrt_ex_1(\prif.rt_ex [1]),
	.prifrt_ex_0(\prif.rt_ex [0]),
	.prifrt_ex_3(\prif.rt_ex [3]),
	.prifrt_ex_2(\prif.rt_ex [2]),
	.prifrt_ex_4(\prif.rt_ex [4]),
	.prifopcode_mem_1(\prif.opcode_mem [1]),
	.prifopcode_mem_0(\prif.opcode_mem [0]),
	.prifopcode_mem_2(\prif.opcode_mem [2]),
	.prifopcode_mem_3(\prif.opcode_mem [3]),
	.prifopcode_mem_5(\prif.opcode_mem [5]),
	.prifopcode_mem_4(\prif.opcode_mem [4]),
	.prifzero_flag_mem(\prif.zero_flag_mem~q ),
	.prifinstr_mem_3(\prif.instr_mem [3]),
	.prifinstr_mem_5(\prif.instr_mem [5]),
	.prifinstr_mem_4(\prif.instr_mem [4]),
	.prifinstr_mem_2(\prif.instr_mem [2]),
	.prifinstr_mem_1(\prif.instr_mem [1]),
	.prifinstr_mem_0(\prif.instr_mem [0]),
	.prifopcode_ex_5(\prif.opcode_ex [5]),
	.prifopcode_ex_0(\prif.opcode_ex [0]),
	.prifopcode_ex_1(\prif.opcode_ex [1]),
	.prifopcode_ex_2(\prif.opcode_ex [2]),
	.prifopcode_ex_4(\prif.opcode_ex [4]),
	.LessThan1(LessThan1),
	.always0(always0),
	.ptBScr(\HU|ptBScr~1_combout ),
	.prifRegwen_wb(\prif.Regwen_wb~q ),
	.prifregwrite_wb_2(\prif.regwrite_wb [2]),
	.prifregwrite_wb_0(\prif.regwrite_wb [0]),
	.prifregwrite_wb_1(\prif.regwrite_wb [1]),
	.prifregwrite_wb_4(\prif.regwrite_wb [4]),
	.prifregwrite_wb_3(\prif.regwrite_wb [3]),
	.Equal8(\HU|Equal8~0_combout ),
	.always01(\HU|always0~5_combout ),
	.prifrs_ex_1(\prif.rs_ex [1]),
	.prifrs_ex_0(\prif.rs_ex [0]),
	.prifrs_ex_3(\prif.rs_ex [3]),
	.prifrs_ex_2(\prif.rs_ex [2]),
	.prifrs_ex_4(\prif.rs_ex [4]),
	.always02(\HU|always0~6_combout ),
	.ptAScr(\HU|ptAScr~4_combout ),
	.always03(always01),
	.exmem_en(\HU|exmem_en~0_combout ),
	.Equal1(\Equal1~1_combout ),
	.ccifiwait_0(ccifiwait_0),
	.always1(\HU|always1~5_combout ),
	.ifid_en(\HU|ifid_en~0_combout ),
	.pc_en(\HU|pc_en~0_combout ),
	.flush_idex(\HU|flush_idex~0_combout ),
	.prifhalt_wb(\prif.halt_wb~q ),
	.ifid_en1(\HU|ifid_en~1_combout ),
	.nRST(nRST),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

pipeline_register PR(
	.prifdmemaddr_1(prifdmemaddr_1),
	.pc_1(pc_1),
	.prifdmemren(prifdmemren),
	.prifdmemwen(prifdmemwen),
	.prifdmemaddr_0(prifdmemaddr_0),
	.pc_0(pc_0),
	.prifdmemaddr_3(prifdmemaddr_3),
	.prifdmemaddr_2(prifdmemaddr_2),
	.prifdmemaddr_5(prifdmemaddr_5),
	.prifdmemaddr_4(prifdmemaddr_4),
	.prifdmemaddr_7(prifdmemaddr_7),
	.prifdmemaddr_6(prifdmemaddr_6),
	.prifdmemaddr_9(prifdmemaddr_9),
	.prifdmemaddr_8(prifdmemaddr_8),
	.prifdmemaddr_11(prifdmemaddr_11),
	.prifdmemaddr_10(prifdmemaddr_10),
	.prifdmemaddr_13(prifdmemaddr_13),
	.prifdmemaddr_12(prifdmemaddr_12),
	.prifdmemaddr_15(prifdmemaddr_15),
	.prifdmemaddr_14(prifdmemaddr_14),
	.prifdmemaddr_23(prifdmemaddr_23),
	.prifdmemaddr_22(prifdmemaddr_22),
	.prifdmemaddr_21(prifdmemaddr_21),
	.prifdmemaddr_29(prifdmemaddr_29),
	.prifdmemaddr_28(prifdmemaddr_28),
	.prifdmemaddr_31(prifdmemaddr_31),
	.prifdmemaddr_30(prifdmemaddr_30),
	.prifdmemaddr_20(prifdmemaddr_20),
	.prifdmemaddr_17(prifdmemaddr_17),
	.prifdmemaddr_16(prifdmemaddr_16),
	.prifdmemaddr_19(prifdmemaddr_19),
	.prifdmemaddr_18(prifdmemaddr_18),
	.prifdmemaddr_25(prifdmemaddr_25),
	.prifdmemaddr_24(prifdmemaddr_24),
	.prifdmemaddr_27(prifdmemaddr_27),
	.prifdmemaddr_26(prifdmemaddr_26),
	.prifhalt_mem(\prif.halt_mem~q ),
	.prifdmemstore_0(prifdmemstore_0),
	.prifimm_ex_1(\prif.imm_ex [1]),
	.prifALUScr_ex_1(\prif.ALUScr_ex [1]),
	.prifshamt_ex_1(\prif.shamt_ex [1]),
	.prifALUScr_ex_0(\prif.ALUScr_ex [0]),
	.prifRegwen_mem(\prif.Regwen_mem~q ),
	.prifregwrite_mem_4(\prif.regwrite_mem [4]),
	.prifregwrite_mem_0(\prif.regwrite_mem [0]),
	.prifregwrite_mem_1(\prif.regwrite_mem [1]),
	.prifregwrite_mem_2(\prif.regwrite_mem [2]),
	.prifregwrite_mem_3(\prif.regwrite_mem [3]),
	.prifrt_ex_1(\prif.rt_ex [1]),
	.prifrt_ex_0(\prif.rt_ex [0]),
	.prifrt_ex_3(\prif.rt_ex [3]),
	.prifrt_ex_2(\prif.rt_ex [2]),
	.prifrt_ex_4(\prif.rt_ex [4]),
	.prifrdat2_ex_1(\prif.rdat2_ex [1]),
	.prifopcode_mem_1(\prif.opcode_mem [1]),
	.prifopcode_mem_0(\prif.opcode_mem [0]),
	.prifopcode_mem_2(\prif.opcode_mem [2]),
	.prifopcode_mem_3(\prif.opcode_mem [3]),
	.prifopcode_mem_5(\prif.opcode_mem [5]),
	.prifopcode_mem_4(\prif.opcode_mem [4]),
	.prifrdat1_ex_1(\prif.rdat1_ex [1]),
	.prifimm_ex_0(\prif.imm_ex [0]),
	.prifshamt_ex_0(\prif.shamt_ex [0]),
	.prifrdat2_ex_0(\prif.rdat2_ex [0]),
	.prifrdat1_ex_0(\prif.rdat1_ex [0]),
	.prifrdat2_ex_3(\prif.rdat2_ex [3]),
	.prifimm_ex_3(\prif.imm_ex [3]),
	.prifshamt_ex_3(\prif.shamt_ex [3]),
	.prifimm_ex_2(\prif.imm_ex [2]),
	.prifshamt_ex_2(\prif.shamt_ex [2]),
	.prifrdat2_ex_2(\prif.rdat2_ex [2]),
	.prifrdat2_ex_4(\prif.rdat2_ex [4]),
	.prifimm_ex_4(\prif.imm_ex [4]),
	.prifshamt_ex_4(\prif.shamt_ex [4]),
	.prifinstr_ex_15(\prif.instr_ex [15]),
	.prifrdat2_ex_31(\prif.rdat2_ex [31]),
	.prifimm_mem_15(\prif.imm_mem [15]),
	.prifrdat2_ex_30(\prif.rdat2_ex [30]),
	.prifimm_mem_14(\prif.imm_mem [14]),
	.prifrdat2_ex_29(\prif.rdat2_ex [29]),
	.prifimm_mem_13(\prif.imm_mem [13]),
	.prifimm_ex_5(\prif.imm_ex [5]),
	.prifrdat2_ex_5(\prif.rdat2_ex [5]),
	.prifimm_ex_15(\prif.imm_ex [15]),
	.prifrdat2_ex_15(\prif.rdat2_ex [15]),
	.prifimm_ex_14(\prif.imm_ex [14]),
	.prifrdat2_ex_14(\prif.rdat2_ex [14]),
	.prifimm_ex_13(\prif.imm_ex [13]),
	.prifrdat2_ex_13(\prif.rdat2_ex [13]),
	.prifimm_ex_12(\prif.imm_ex [12]),
	.prifrdat2_ex_12(\prif.rdat2_ex [12]),
	.prifimm_ex_11(\prif.imm_ex [11]),
	.prifrdat2_ex_11(\prif.rdat2_ex [11]),
	.prifimm_ex_10(\prif.imm_ex [10]),
	.prifrdat2_ex_10(\prif.rdat2_ex [10]),
	.prifimm_ex_9(\prif.imm_ex [9]),
	.prifrdat2_ex_9(\prif.rdat2_ex [9]),
	.prifimm_ex_6(\prif.imm_ex [6]),
	.prifrdat2_ex_6(\prif.rdat2_ex [6]),
	.prifrdat2_ex_27(\prif.rdat2_ex [27]),
	.prifimm_mem_11(\prif.imm_mem [11]),
	.prifrdat2_ex_23(\prif.rdat2_ex [23]),
	.prifimm_mem_7(\prif.imm_mem [7]),
	.prifrdat2_ex_18(\prif.rdat2_ex [18]),
	.prifimm_mem_2(\prif.imm_mem [2]),
	.prifrdat2_ex_24(\prif.rdat2_ex [24]),
	.prifimm_mem_8(\prif.imm_mem [8]),
	.prifrdat2_ex_16(\prif.rdat2_ex [16]),
	.prifimm_mem_0(\prif.imm_mem [0]),
	.prifrdat2_ex_19(\prif.rdat2_ex [19]),
	.prifimm_mem_3(\prif.imm_mem [3]),
	.prifrdat2_ex_17(\prif.rdat2_ex [17]),
	.prifimm_mem_1(\prif.imm_mem [1]),
	.prifrdat2_ex_21(\prif.rdat2_ex [21]),
	.prifimm_mem_5(\prif.imm_mem [5]),
	.prifrdat2_ex_20(\prif.rdat2_ex [20]),
	.prifimm_mem_4(\prif.imm_mem [4]),
	.prifrdat2_ex_28(\prif.rdat2_ex [28]),
	.prifimm_mem_12(\prif.imm_mem [12]),
	.prifrdat2_ex_26(\prif.rdat2_ex [26]),
	.prifimm_mem_10(\prif.imm_mem [10]),
	.prifimm_ex_8(\prif.imm_ex [8]),
	.prifrdat2_ex_8(\prif.rdat2_ex [8]),
	.prifimm_ex_7(\prif.imm_ex [7]),
	.prifrdat2_ex_7(\prif.rdat2_ex [7]),
	.prifrdat2_ex_22(\prif.rdat2_ex [22]),
	.prifimm_mem_6(\prif.imm_mem [6]),
	.prifrdat2_ex_25(\prif.rdat2_ex [25]),
	.prifimm_mem_9(\prif.imm_mem [9]),
	.prifrdat1_ex_2(\prif.rdat1_ex [2]),
	.prifrdat1_ex_4(\prif.rdat1_ex [4]),
	.prifrdat1_ex_3(\prif.rdat1_ex [3]),
	.prifrdat1_ex_8(\prif.rdat1_ex [8]),
	.prifrdat1_ex_7(\prif.rdat1_ex [7]),
	.prifrdat1_ex_6(\prif.rdat1_ex [6]),
	.prifrdat1_ex_5(\prif.rdat1_ex [5]),
	.prifrdat1_ex_16(\prif.rdat1_ex [16]),
	.prifrdat1_ex_15(\prif.rdat1_ex [15]),
	.prifrdat1_ex_14(\prif.rdat1_ex [14]),
	.prifrdat1_ex_13(\prif.rdat1_ex [13]),
	.prifrdat1_ex_11(\prif.rdat1_ex [11]),
	.prifrdat1_ex_12(\prif.rdat1_ex [12]),
	.prifrdat1_ex_10(\prif.rdat1_ex [10]),
	.prifrdat1_ex_9(\prif.rdat1_ex [9]),
	.prifrdat1_ex_18(\prif.rdat1_ex [18]),
	.prifrdat1_ex_17(\prif.rdat1_ex [17]),
	.prifrdat1_ex_20(\prif.rdat1_ex [20]),
	.prifrdat1_ex_19(\prif.rdat1_ex [19]),
	.prifrdat1_ex_22(\prif.rdat1_ex [22]),
	.prifrdat1_ex_21(\prif.rdat1_ex [21]),
	.prifrdat1_ex_24(\prif.rdat1_ex [24]),
	.prifrdat1_ex_23(\prif.rdat1_ex [23]),
	.prifrdat1_ex_31(\prif.rdat1_ex [31]),
	.prifrdat1_ex_30(\prif.rdat1_ex [30]),
	.prifrdat1_ex_29(\prif.rdat1_ex [29]),
	.prifrdat1_ex_26(\prif.rdat1_ex [26]),
	.prifrdat1_ex_25(\prif.rdat1_ex [25]),
	.prifrdat1_ex_28(\prif.rdat1_ex [28]),
	.prifrdat1_ex_27(\prif.rdat1_ex [27]),
	.prifzero_flag_mem(\prif.zero_flag_mem~q ),
	.prifinstr_mem_3(\prif.instr_mem [3]),
	.prifinstr_mem_5(\prif.instr_mem [5]),
	.prifinstr_mem_4(\prif.instr_mem [4]),
	.prifinstr_mem_2(\prif.instr_mem [2]),
	.prifinstr_mem_1(\prif.instr_mem [1]),
	.prifinstr_mem_0(\prif.instr_mem [0]),
	.prifrdat1_mem_1(\prif.rdat1_mem [1]),
	.prifPCScr_mem_0(\prif.PCScr_mem [0]),
	.prifpc_bran_mem_1(\prif.pc_bran_mem [1]),
	.prifPCScr_mem_1(\prif.PCScr_mem [1]),
	.prifopcode_ex_5(\prif.opcode_ex [5]),
	.prifopcode_ex_0(\prif.opcode_ex [0]),
	.prifopcode_ex_1(\prif.opcode_ex [1]),
	.prifopcode_ex_2(\prif.opcode_ex [2]),
	.prifopcode_ex_4(\prif.opcode_ex [4]),
	.prifmemren_ex(\prif.memren_ex~q ),
	.prifmemwen_ex(\prif.memwen_ex~q ),
	.prifrdat1_mem_0(\prif.rdat1_mem [0]),
	.prifpc_bran_mem_0(\prif.pc_bran_mem [0]),
	.prifrdat1_mem_3(\prif.rdat1_mem [3]),
	.prifpc_bran_mem_3(\prif.pc_bran_mem [3]),
	.prifrdat1_mem_2(\prif.rdat1_mem [2]),
	.prifpc_bran_mem_2(\prif.pc_bran_mem [2]),
	.prifrdat1_mem_5(\prif.rdat1_mem [5]),
	.prifpc_bran_mem_5(\prif.pc_bran_mem [5]),
	.prifrdat1_mem_4(\prif.rdat1_mem [4]),
	.prifpc_bran_mem_4(\prif.pc_bran_mem [4]),
	.prifrdat1_mem_7(\prif.rdat1_mem [7]),
	.prifpc_bran_mem_7(\prif.pc_bran_mem [7]),
	.prifrdat1_mem_6(\prif.rdat1_mem [6]),
	.prifpc_bran_mem_6(\prif.pc_bran_mem [6]),
	.prifrdat1_mem_9(\prif.rdat1_mem [9]),
	.prifpc_bran_mem_9(\prif.pc_bran_mem [9]),
	.prifinstr_mem_7(\prif.instr_mem [7]),
	.prifrdat1_mem_8(\prif.rdat1_mem [8]),
	.prifpc_bran_mem_8(\prif.pc_bran_mem [8]),
	.prifinstr_mem_6(\prif.instr_mem [6]),
	.prifrdat1_mem_11(\prif.rdat1_mem [11]),
	.prifpc_bran_mem_11(\prif.pc_bran_mem [11]),
	.prifinstr_mem_9(\prif.instr_mem [9]),
	.prifrdat1_mem_10(\prif.rdat1_mem [10]),
	.prifpc_bran_mem_10(\prif.pc_bran_mem [10]),
	.prifinstr_mem_8(\prif.instr_mem [8]),
	.prifrdat1_mem_13(\prif.rdat1_mem [13]),
	.prifpc_bran_mem_13(\prif.pc_bran_mem [13]),
	.prifinstr_mem_11(\prif.instr_mem [11]),
	.prifrdat1_mem_12(\prif.rdat1_mem [12]),
	.prifpc_bran_mem_12(\prif.pc_bran_mem [12]),
	.prifinstr_mem_10(\prif.instr_mem [10]),
	.prifrdat1_mem_15(\prif.rdat1_mem [15]),
	.prifpc_bran_mem_15(\prif.pc_bran_mem [15]),
	.prifinstr_mem_13(\prif.instr_mem [13]),
	.prifrdat1_mem_14(\prif.rdat1_mem [14]),
	.prifpc_bran_mem_14(\prif.pc_bran_mem [14]),
	.prifinstr_mem_12(\prif.instr_mem [12]),
	.prifrdat1_mem_23(\prif.rdat1_mem [23]),
	.prifpc_bran_mem_23(\prif.pc_bran_mem [23]),
	.prifinstr_mem_21(\prif.instr_mem [21]),
	.prifrdat1_mem_22(\prif.rdat1_mem [22]),
	.prifpc_bran_mem_22(\prif.pc_bran_mem [22]),
	.prifinstr_mem_20(\prif.instr_mem [20]),
	.prifrdat1_mem_21(\prif.rdat1_mem [21]),
	.prifpc_bran_mem_21(\prif.pc_bran_mem [21]),
	.prifinstr_mem_19(\prif.instr_mem [19]),
	.prifrdat1_mem_29(\prif.rdat1_mem [29]),
	.prifpc_bran_mem_29(\prif.pc_bran_mem [29]),
	.prifrdat1_mem_28(\prif.rdat1_mem [28]),
	.prifpc_bran_mem_28(\prif.pc_bran_mem [28]),
	.prifrdat1_mem_31(\prif.rdat1_mem [31]),
	.prifpc_bran_mem_31(\prif.pc_bran_mem [31]),
	.prifrdat1_mem_30(\prif.rdat1_mem [30]),
	.prifpc_bran_mem_30(\prif.pc_bran_mem [30]),
	.prifrdat1_mem_20(\prif.rdat1_mem [20]),
	.prifpc_bran_mem_20(\prif.pc_bran_mem [20]),
	.prifinstr_mem_18(\prif.instr_mem [18]),
	.prifrdat1_mem_17(\prif.rdat1_mem [17]),
	.prifpc_bran_mem_17(\prif.pc_bran_mem [17]),
	.prifinstr_mem_15(\prif.instr_mem [15]),
	.prifrdat1_mem_16(\prif.rdat1_mem [16]),
	.prifpc_bran_mem_16(\prif.pc_bran_mem [16]),
	.prifinstr_mem_14(\prif.instr_mem [14]),
	.prifrdat1_mem_19(\prif.rdat1_mem [19]),
	.prifpc_bran_mem_19(\prif.pc_bran_mem [19]),
	.prifinstr_mem_17(\prif.instr_mem [17]),
	.prifrdat1_mem_18(\prif.rdat1_mem [18]),
	.prifpc_bran_mem_18(\prif.pc_bran_mem [18]),
	.prifinstr_mem_16(\prif.instr_mem [16]),
	.prifrdat1_mem_25(\prif.rdat1_mem [25]),
	.prifpc_bran_mem_25(\prif.pc_bran_mem [25]),
	.prifinstr_mem_23(\prif.instr_mem [23]),
	.prifrdat1_mem_24(\prif.rdat1_mem [24]),
	.prifpc_bran_mem_24(\prif.pc_bran_mem [24]),
	.prifinstr_mem_22(\prif.instr_mem [22]),
	.prifrdat1_mem_27(\prif.rdat1_mem [27]),
	.prifpc_bran_mem_27(\prif.pc_bran_mem [27]),
	.prifinstr_mem_25(\prif.instr_mem [25]),
	.prifrdat1_mem_26(\prif.rdat1_mem [26]),
	.prifpc_bran_mem_26(\prif.pc_bran_mem [26]),
	.prifinstr_mem_24(\prif.instr_mem [24]),
	.prifdmemstore_1(prifdmemstore_1),
	.prifdmemstore_2(prifdmemstore_2),
	.prifdmemstore_3(prifdmemstore_3),
	.prifdmemstore_4(prifdmemstore_4),
	.prifdmemstore_5(prifdmemstore_5),
	.prifdmemstore_6(prifdmemstore_6),
	.prifdmemstore_7(prifdmemstore_7),
	.prifdmemstore_8(prifdmemstore_8),
	.prifdmemstore_9(prifdmemstore_9),
	.prifdmemstore_10(prifdmemstore_10),
	.prifdmemstore_11(prifdmemstore_11),
	.prifdmemstore_12(prifdmemstore_12),
	.prifdmemstore_13(prifdmemstore_13),
	.prifdmemstore_14(prifdmemstore_14),
	.prifdmemstore_15(prifdmemstore_15),
	.prifdmemstore_16(prifdmemstore_16),
	.prifdmemstore_17(prifdmemstore_17),
	.prifdmemstore_18(prifdmemstore_18),
	.prifdmemstore_19(prifdmemstore_19),
	.prifdmemstore_20(prifdmemstore_20),
	.prifdmemstore_21(prifdmemstore_21),
	.prifdmemstore_22(prifdmemstore_22),
	.prifdmemstore_23(prifdmemstore_23),
	.prifdmemstore_24(prifdmemstore_24),
	.prifdmemstore_25(prifdmemstore_25),
	.prifdmemstore_26(prifdmemstore_26),
	.prifdmemstore_27(prifdmemstore_27),
	.prifdmemstore_28(prifdmemstore_28),
	.prifdmemstore_29(prifdmemstore_29),
	.prifdmemstore_30(prifdmemstore_30),
	.prifdmemstore_31(prifdmemstore_31),
	.prifhalt_ex(\prif.halt_ex~q ),
	.prifimemload_id_31(\prif.imemload_id [31]),
	.prifimemload_id_30(\prif.imemload_id [30]),
	.prifimemload_id_29(\prif.imemload_id [29]),
	.prifimemload_id_27(\prif.imemload_id [27]),
	.prifimemload_id_26(\prif.imemload_id [26]),
	.prifimemload_id_28(\prif.imemload_id [28]),
	.prifimemload_id_3(\prif.imemload_id [3]),
	.prifimemload_id_1(\prif.imemload_id [1]),
	.prifimemload_id_5(\prif.imemload_id [5]),
	.prifimemload_id_4(\prif.imemload_id [4]),
	.prifimemload_id_2(\prif.imemload_id [2]),
	.prifimemload_id_0(\prif.imemload_id [0]),
	.prifimemload_id_7(\prif.imemload_id [7]),
	.prifRegwen_ex(\prif.Regwen_ex~q ),
	.prifrd_ex_4(\prif.rd_ex [4]),
	.prifRegDest_ex_1(\prif.RegDest_ex [1]),
	.prifRegDest_ex_0(\prif.RegDest_ex [0]),
	.prifrd_ex_0(\prif.rd_ex [0]),
	.prifrd_ex_1(\prif.rd_ex [1]),
	.prifrd_ex_2(\prif.rd_ex [2]),
	.prifrd_ex_3(\prif.rd_ex [3]),
	.prifimemload_id_17(\prif.imemload_id [17]),
	.prifimemload_id_16(\prif.imemload_id [16]),
	.prifimemload_id_19(\prif.imemload_id [19]),
	.prifimemload_id_18(\prif.imemload_id [18]),
	.prifimemload_id_20(\prif.imemload_id [20]),
	.prifdataScr_mem_0(\prif.dataScr_mem [0]),
	.prifdataScr_mem_1(\prif.dataScr_mem [1]),
	.prifimemload_id_22(\prif.imemload_id [22]),
	.prifimemload_id_21(\prif.imemload_id [21]),
	.prifimemload_id_24(\prif.imemload_id [24]),
	.prifimemload_id_23(\prif.imemload_id [23]),
	.prifimemload_id_25(\prif.imemload_id [25]),
	.prifopcode_ex_3(\prif.opcode_ex [3]),
	.prifimemload_id_6(\prif.imemload_id [6]),
	.prifimemload_id_9(\prif.imemload_id [9]),
	.prifimemload_id_8(\prif.imemload_id [8]),
	.prifimemload_id_10(\prif.imemload_id [10]),
	.prifimemload_id_15(\prif.imemload_id [15]),
	.prifimemload_id_14(\prif.imemload_id [14]),
	.prifimemload_id_13(\prif.imemload_id [13]),
	.prifimemload_id_12(\prif.imemload_id [12]),
	.prifimemload_id_11(\prif.imemload_id [11]),
	.prifinstr_ex_3(\prif.instr_ex [3]),
	.prifinstr_ex_5(\prif.instr_ex [5]),
	.prifinstr_ex_4(\prif.instr_ex [4]),
	.prifinstr_ex_2(\prif.instr_ex [2]),
	.prifinstr_ex_1(\prif.instr_ex [1]),
	.prifinstr_ex_0(\prif.instr_ex [0]),
	.prifPCScr_ex_0(\prif.PCScr_ex [0]),
	.prifpc_ex_1(\prif.pc_ex [1]),
	.prifPCScr_ex_1(\prif.PCScr_ex [1]),
	.prifpc_ex_0(\prif.pc_ex [0]),
	.prifpc_ex_3(\prif.pc_ex [3]),
	.prifpc_ex_2(\prif.pc_ex [2]),
	.Add0(\Add0~0_combout ),
	.Add01(\Add0~2_combout ),
	.prifpc_ex_5(\prif.pc_ex [5]),
	.prifpc_ex_4(\prif.pc_ex [4]),
	.Add02(\Add0~4_combout ),
	.Add03(\Add0~6_combout ),
	.prifpc_ex_7(\prif.pc_ex [7]),
	.prifpc_ex_6(\prif.pc_ex [6]),
	.Add04(\Add0~8_combout ),
	.Add05(\Add0~10_combout ),
	.prifpc_ex_9(\prif.pc_ex [9]),
	.prifpc_ex_8(\prif.pc_ex [8]),
	.Add06(\Add0~12_combout ),
	.Add07(\Add0~14_combout ),
	.prifinstr_ex_7(\prif.instr_ex [7]),
	.prifinstr_ex_6(\prif.instr_ex [6]),
	.prifpc_ex_11(\prif.pc_ex [11]),
	.prifpc_ex_10(\prif.pc_ex [10]),
	.Add08(\Add0~16_combout ),
	.Add09(\Add0~18_combout ),
	.prifinstr_ex_9(\prif.instr_ex [9]),
	.prifinstr_ex_8(\prif.instr_ex [8]),
	.prifpc_ex_13(\prif.pc_ex [13]),
	.prifpc_ex_12(\prif.pc_ex [12]),
	.Add010(\Add0~20_combout ),
	.Add011(\Add0~22_combout ),
	.prifinstr_ex_11(\prif.instr_ex [11]),
	.prifinstr_ex_10(\prif.instr_ex [10]),
	.prifpc_ex_15(\prif.pc_ex [15]),
	.prifpc_ex_14(\prif.pc_ex [14]),
	.Add012(\Add0~24_combout ),
	.Add013(\Add0~26_combout ),
	.prifinstr_ex_13(\prif.instr_ex [13]),
	.prifinstr_ex_12(\prif.instr_ex [12]),
	.prifpc_ex_23(\prif.pc_ex [23]),
	.prifpc_ex_22(\prif.pc_ex [22]),
	.prifpc_ex_21(\prif.pc_ex [21]),
	.prifpc_ex_20(\prif.pc_ex [20]),
	.prifpc_ex_19(\prif.pc_ex [19]),
	.prifpc_ex_18(\prif.pc_ex [18]),
	.prifpc_ex_17(\prif.pc_ex [17]),
	.prifpc_ex_16(\prif.pc_ex [16]),
	.Add014(\Add0~28_combout ),
	.Add015(\Add0~30_combout ),
	.Add016(\Add0~32_combout ),
	.Add017(\Add0~34_combout ),
	.Add018(\Add0~36_combout ),
	.Add019(\Add0~38_combout ),
	.Add020(\Add0~40_combout ),
	.Add021(\Add0~42_combout ),
	.prifinstr_ex_21(\prif.instr_ex [21]),
	.prifinstr_ex_20(\prif.instr_ex [20]),
	.prifinstr_ex_19(\prif.instr_ex [19]),
	.prifpc_ex_29(\prif.pc_ex [29]),
	.prifpc_ex_28(\prif.pc_ex [28]),
	.prifpc_ex_27(\prif.pc_ex [27]),
	.prifpc_ex_26(\prif.pc_ex [26]),
	.prifpc_ex_25(\prif.pc_ex [25]),
	.prifpc_ex_24(\prif.pc_ex [24]),
	.Add022(\Add0~44_combout ),
	.Add023(\Add0~46_combout ),
	.Add024(\Add0~48_combout ),
	.Add025(\Add0~50_combout ),
	.Add026(\Add0~52_combout ),
	.Add027(\Add0~54_combout ),
	.prifpc_ex_31(\prif.pc_ex [31]),
	.prifpc_ex_30(\prif.pc_ex [30]),
	.Add028(\Add0~56_combout ),
	.Add029(\Add0~58_combout ),
	.prifinstr_ex_18(\prif.instr_ex [18]),
	.prifinstr_ex_14(\prif.instr_ex [14]),
	.prifinstr_ex_17(\prif.instr_ex [17]),
	.prifinstr_ex_16(\prif.instr_ex [16]),
	.prifinstr_ex_23(\prif.instr_ex [23]),
	.prifinstr_ex_22(\prif.instr_ex [22]),
	.prifinstr_ex_25(\prif.instr_ex [25]),
	.prifinstr_ex_24(\prif.instr_ex [24]),
	.prifdataScr_ex_0(\prif.dataScr_ex [0]),
	.prifdataScr_ex_1(\prif.dataScr_ex [1]),
	.prifpc_id_1(\prif.pc_id [1]),
	.prifpc_id_0(\prif.pc_id [0]),
	.prifpc_id_3(\prif.pc_id [3]),
	.prifpc_id_2(\prif.pc_id [2]),
	.prifpc_id_5(\prif.pc_id [5]),
	.prifpc_id_4(\prif.pc_id [4]),
	.prifpc_id_7(\prif.pc_id [7]),
	.prifpc_id_6(\prif.pc_id [6]),
	.prifpc_id_9(\prif.pc_id [9]),
	.prifpc_id_8(\prif.pc_id [8]),
	.prifpc_id_11(\prif.pc_id [11]),
	.prifpc_id_10(\prif.pc_id [10]),
	.prifpc_id_13(\prif.pc_id [13]),
	.prifpc_id_12(\prif.pc_id [12]),
	.prifpc_id_15(\prif.pc_id [15]),
	.prifpc_id_14(\prif.pc_id [14]),
	.prifpc_id_23(\prif.pc_id [23]),
	.prifpc_id_22(\prif.pc_id [22]),
	.prifpc_id_21(\prif.pc_id [21]),
	.prifpc_id_20(\prif.pc_id [20]),
	.prifpc_id_19(\prif.pc_id [19]),
	.prifpc_id_18(\prif.pc_id [18]),
	.prifpc_id_17(\prif.pc_id [17]),
	.prifpc_id_16(\prif.pc_id [16]),
	.prifpc_id_29(\prif.pc_id [29]),
	.prifpc_id_28(\prif.pc_id [28]),
	.prifpc_id_27(\prif.pc_id [27]),
	.prifpc_id_26(\prif.pc_id [26]),
	.prifpc_id_25(\prif.pc_id [25]),
	.prifpc_id_24(\prif.pc_id [24]),
	.prifpc_id_31(\prif.pc_id [31]),
	.prifpc_id_30(\prif.pc_id [30]),
	.Add2(\Add2~0_combout ),
	.Add21(\Add2~2_combout ),
	.Add22(\Add2~4_combout ),
	.Add23(\Add2~6_combout ),
	.Add24(\Add2~8_combout ),
	.Add25(\Add2~10_combout ),
	.Add26(\Add2~12_combout ),
	.Add27(\Add2~14_combout ),
	.Add28(\Add2~16_combout ),
	.Add29(\Add2~18_combout ),
	.Add210(\Add2~20_combout ),
	.Add211(\Add2~22_combout ),
	.Add212(\Add2~24_combout ),
	.Add213(\Add2~26_combout ),
	.Add214(\Add2~28_combout ),
	.Add215(\Add2~30_combout ),
	.Add216(\Add2~32_combout ),
	.Add217(\Add2~34_combout ),
	.Add218(\Add2~36_combout ),
	.Add219(\Add2~38_combout ),
	.Add220(\Add2~40_combout ),
	.Add221(\Add2~42_combout ),
	.Add222(\Add2~44_combout ),
	.Add223(\Add2~46_combout ),
	.Add224(\Add2~48_combout ),
	.Add225(\Add2~50_combout ),
	.Add226(\Add2~52_combout ),
	.Add227(\Add2~54_combout ),
	.Add228(\Add2~56_combout ),
	.pc_2(pc_2),
	.always1(always1),
	.ramiframload_0(ramiframload_0),
	.ramiframload_1(ramiframload_1),
	.ramiframload_2(ramiframload_2),
	.ramiframload_3(ramiframload_3),
	.ramiframload_4(ramiframload_4),
	.ramiframload_5(ramiframload_5),
	.ramiframload_6(ramiframload_6),
	.ramiframload_7(ramiframload_7),
	.ramiframload_8(ramiframload_8),
	.ramiframload_9(ramiframload_9),
	.ramiframload_10(ramiframload_10),
	.ramiframload_11(ramiframload_11),
	.ramiframload_12(ramiframload_12),
	.ramiframload_13(ramiframload_13),
	.ramiframload_14(ramiframload_14),
	.ramiframload_15(ramiframload_15),
	.ramiframload_16(ramiframload_16),
	.ramiframload_17(ramiframload_17),
	.ramiframload_18(ramiframload_18),
	.ramiframload_19(ramiframload_19),
	.ramiframload_20(ramiframload_20),
	.ramiframload_21(ramiframload_21),
	.ramiframload_22(ramiframload_22),
	.ramiframload_23(ramiframload_23),
	.ramiframload_24(ramiframload_24),
	.ramiframload_25(ramiframload_25),
	.ramiframload_26(ramiframload_26),
	.ramiframload_27(ramiframload_27),
	.ramiframload_28(ramiframload_28),
	.ramiframload_29(ramiframload_29),
	.ramiframload_30(ramiframload_30),
	.ramiframload_31(ramiframload_31),
	.prifALUOP_ex_3(\prif.ALUOP_ex [3]),
	.prifRegwen_wb(\prif.Regwen_wb~q ),
	.prifregwrite_wb_2(\prif.regwrite_wb [2]),
	.prifregwrite_wb_0(\prif.regwrite_wb [0]),
	.prifregwrite_wb_1(\prif.regwrite_wb [1]),
	.prifregwrite_wb_4(\prif.regwrite_wb [4]),
	.prifregwrite_wb_3(\prif.regwrite_wb [3]),
	.Mux62(\Mux62~0_combout ),
	.prifdmemload_wb_1(\prif.dmemload_wb [1]),
	.prifdmemaddr_wb_1(\prif.dmemaddr_wb [1]),
	.prifdataScr_wb_0(\prif.dataScr_wb [0]),
	.prifdataScr_wb_1(\prif.dataScr_wb [1]),
	.prifpc_wb_1(\prif.pc_wb [1]),
	.Mux621(\Mux62~1_combout ),
	.prifrs_ex_1(\prif.rs_ex [1]),
	.prifrs_ex_0(\prif.rs_ex [0]),
	.prifrs_ex_3(\prif.rs_ex [3]),
	.prifrs_ex_2(\prif.rs_ex [2]),
	.prifrs_ex_4(\prif.rs_ex [4]),
	.Mux63(\Mux63~0_combout ),
	.prifdmemload_wb_0(\prif.dmemload_wb [0]),
	.prifdmemaddr_wb_0(\prif.dmemaddr_wb [0]),
	.prifpc_wb_0(\prif.pc_wb [0]),
	.Mux631(\Mux63~1_combout ),
	.prifdmemload_wb_3(\prif.dmemload_wb [3]),
	.prifdmemaddr_wb_3(\prif.dmemaddr_wb [3]),
	.prifpc_wb_3(\prif.pc_wb [3]),
	.prifdmemload_wb_2(\prif.dmemload_wb [2]),
	.prifdmemaddr_wb_2(\prif.dmemaddr_wb [2]),
	.prifpc_wb_2(\prif.pc_wb [2]),
	.Mux61(\Mux61~1_combout ),
	.prifdmemload_wb_4(\prif.dmemload_wb [4]),
	.prifdmemaddr_wb_4(\prif.dmemaddr_wb [4]),
	.prifpc_wb_4(\prif.pc_wb [4]),
	.prifdmemload_wb_31(\prif.dmemload_wb [31]),
	.prifimm_wb_15(\prif.imm_wb [15]),
	.prifdmemaddr_wb_31(\prif.dmemaddr_wb [31]),
	.prifpc_wb_31(\prif.pc_wb [31]),
	.Mux32(\Mux32~1_combout ),
	.prifimm_wb_14(\prif.imm_wb [14]),
	.prifdmemload_wb_30(\prif.dmemload_wb [30]),
	.prifdmemaddr_wb_30(\prif.dmemaddr_wb [30]),
	.prifpc_wb_30(\prif.pc_wb [30]),
	.Mux33(\Mux33~1_combout ),
	.prifdmemload_wb_29(\prif.dmemload_wb [29]),
	.prifimm_wb_13(\prif.imm_wb [13]),
	.prifdmemaddr_wb_29(\prif.dmemaddr_wb [29]),
	.prifpc_wb_29(\prif.pc_wb [29]),
	.Mux34(\Mux34~1_combout ),
	.prifdmemload_wb_5(\prif.dmemload_wb [5]),
	.prifdmemaddr_wb_5(\prif.dmemaddr_wb [5]),
	.prifpc_wb_5(\prif.pc_wb [5]),
	.prifdmemload_wb_15(\prif.dmemload_wb [15]),
	.prifdmemaddr_wb_15(\prif.dmemaddr_wb [15]),
	.prifpc_wb_15(\prif.pc_wb [15]),
	.prifdmemload_wb_14(\prif.dmemload_wb [14]),
	.prifdmemaddr_wb_14(\prif.dmemaddr_wb [14]),
	.prifpc_wb_14(\prif.pc_wb [14]),
	.prifdmemload_wb_13(\prif.dmemload_wb [13]),
	.prifdmemaddr_wb_13(\prif.dmemaddr_wb [13]),
	.prifpc_wb_13(\prif.pc_wb [13]),
	.prifdmemload_wb_12(\prif.dmemload_wb [12]),
	.prifdmemaddr_wb_12(\prif.dmemaddr_wb [12]),
	.prifpc_wb_12(\prif.pc_wb [12]),
	.prifdmemload_wb_11(\prif.dmemload_wb [11]),
	.prifdmemaddr_wb_11(\prif.dmemaddr_wb [11]),
	.prifpc_wb_11(\prif.pc_wb [11]),
	.prifdmemload_wb_10(\prif.dmemload_wb [10]),
	.prifdmemaddr_wb_10(\prif.dmemaddr_wb [10]),
	.prifpc_wb_10(\prif.pc_wb [10]),
	.prifdmemload_wb_9(\prif.dmemload_wb [9]),
	.prifdmemaddr_wb_9(\prif.dmemaddr_wb [9]),
	.prifpc_wb_9(\prif.pc_wb [9]),
	.prifdmemload_wb_6(\prif.dmemload_wb [6]),
	.prifdmemaddr_wb_6(\prif.dmemaddr_wb [6]),
	.prifpc_wb_6(\prif.pc_wb [6]),
	.prifdmemload_wb_27(\prif.dmemload_wb [27]),
	.prifimm_wb_11(\prif.imm_wb [11]),
	.prifdmemaddr_wb_27(\prif.dmemaddr_wb [27]),
	.prifpc_wb_27(\prif.pc_wb [27]),
	.Mux36(\Mux36~1_combout ),
	.prifdmemload_wb_23(\prif.dmemload_wb [23]),
	.prifimm_wb_7(\prif.imm_wb [7]),
	.prifdmemaddr_wb_23(\prif.dmemaddr_wb [23]),
	.prifpc_wb_23(\prif.pc_wb [23]),
	.Mux40(\Mux40~1_combout ),
	.prifimm_wb_2(\prif.imm_wb [2]),
	.prifdmemload_wb_18(\prif.dmemload_wb [18]),
	.prifdmemaddr_wb_18(\prif.dmemaddr_wb [18]),
	.prifpc_wb_18(\prif.pc_wb [18]),
	.Mux45(\Mux45~1_combout ),
	.prifimm_wb_8(\prif.imm_wb [8]),
	.prifdmemload_wb_24(\prif.dmemload_wb [24]),
	.prifdmemaddr_wb_24(\prif.dmemaddr_wb [24]),
	.prifpc_wb_24(\prif.pc_wb [24]),
	.Mux39(\Mux39~1_combout ),
	.prifimm_wb_0(\prif.imm_wb [0]),
	.prifdmemload_wb_16(\prif.dmemload_wb [16]),
	.prifdmemaddr_wb_16(\prif.dmemaddr_wb [16]),
	.prifpc_wb_16(\prif.pc_wb [16]),
	.Mux47(\Mux47~1_combout ),
	.prifdmemload_wb_19(\prif.dmemload_wb [19]),
	.prifimm_wb_3(\prif.imm_wb [3]),
	.prifdmemaddr_wb_19(\prif.dmemaddr_wb [19]),
	.prifpc_wb_19(\prif.pc_wb [19]),
	.Mux44(\Mux44~1_combout ),
	.prifdmemload_wb_17(\prif.dmemload_wb [17]),
	.prifimm_wb_1(\prif.imm_wb [1]),
	.prifdmemaddr_wb_17(\prif.dmemaddr_wb [17]),
	.prifpc_wb_17(\prif.pc_wb [17]),
	.Mux46(\Mux46~1_combout ),
	.prifdmemload_wb_21(\prif.dmemload_wb [21]),
	.prifimm_wb_5(\prif.imm_wb [5]),
	.prifdmemaddr_wb_21(\prif.dmemaddr_wb [21]),
	.prifpc_wb_21(\prif.pc_wb [21]),
	.Mux42(\Mux42~1_combout ),
	.prifimm_wb_4(\prif.imm_wb [4]),
	.prifdmemload_wb_20(\prif.dmemload_wb [20]),
	.prifdmemaddr_wb_20(\prif.dmemaddr_wb [20]),
	.prifpc_wb_20(\prif.pc_wb [20]),
	.Mux43(\Mux43~1_combout ),
	.prifimm_wb_12(\prif.imm_wb [12]),
	.prifdmemload_wb_28(\prif.dmemload_wb [28]),
	.prifdmemaddr_wb_28(\prif.dmemaddr_wb [28]),
	.prifpc_wb_28(\prif.pc_wb [28]),
	.Mux35(\Mux35~1_combout ),
	.prifimm_wb_10(\prif.imm_wb [10]),
	.prifdmemload_wb_26(\prif.dmemload_wb [26]),
	.prifdmemaddr_wb_26(\prif.dmemaddr_wb [26]),
	.prifpc_wb_26(\prif.pc_wb [26]),
	.Mux37(\Mux37~1_combout ),
	.prifdmemload_wb_8(\prif.dmemload_wb [8]),
	.prifdmemaddr_wb_8(\prif.dmemaddr_wb [8]),
	.prifpc_wb_8(\prif.pc_wb [8]),
	.prifdmemload_wb_7(\prif.dmemload_wb [7]),
	.prifdmemaddr_wb_7(\prif.dmemaddr_wb [7]),
	.prifpc_wb_7(\prif.pc_wb [7]),
	.prifimm_wb_6(\prif.imm_wb [6]),
	.prifdmemload_wb_22(\prif.dmemload_wb [22]),
	.prifdmemaddr_wb_22(\prif.dmemaddr_wb [22]),
	.prifpc_wb_22(\prif.pc_wb [22]),
	.Mux41(\Mux41~1_combout ),
	.prifdmemload_wb_25(\prif.dmemload_wb [25]),
	.prifimm_wb_9(\prif.imm_wb [9]),
	.prifdmemaddr_wb_25(\prif.dmemaddr_wb [25]),
	.prifpc_wb_25(\prif.pc_wb [25]),
	.Mux38(\Mux38~1_combout ),
	.prifALUOP_ex_2(\prif.ALUOP_ex [2]),
	.prifALUOP_ex_1(\prif.ALUOP_ex [1]),
	.prifALUOP_ex_0(\prif.ALUOP_ex [0]),
	.aluifportOut_1(\ALU|aluif.portOut[1]~15_combout ),
	.exmem_en(\HU|exmem_en~0_combout ),
	.dmemaddr(\PR|dmemaddr~0_combout ),
	.ccifiwait_0(ccifiwait_0),
	.dmemren(\PR|dmemren~0_combout ),
	.dmemwen(\PR|dmemwen~0_combout ),
	.aluifportOut_0(\ALU|aluif.portOut[0]~24_combout ),
	.dmemaddr1(\PR|dmemaddr~1_combout ),
	.aluifportOut_3(\ALU|aluif.portOut[3]~30_combout ),
	.aluifportOut_5(\ALU|aluif.portOut[5]~31_combout ),
	.aluifportOut_2(\ALU|aluif.portOut[2]~33_combout ),
	.aluifportOut_31(\ALU|aluif.portOut[3]~39_combout ),
	.aluifportOut_32(\ALU|aluif.portOut[3]~40_combout ),
	.dmemaddr2(\PR|dmemaddr~2_combout ),
	.aluifportOut_21(\ALU|aluif.portOut[2]~48_combout ),
	.dmemaddr3(\PR|dmemaddr~3_combout ),
	.aluifportOut_51(\ALU|aluif.portOut[5]~57_combout ),
	.aluifportOut_52(\ALU|aluif.portOut[5]~58_combout ),
	.dmemaddr4(\PR|dmemaddr~4_combout ),
	.aluifportOut_4(\ALU|aluif.portOut[4]~65_combout ),
	.dmemaddr5(\PR|dmemaddr~5_combout ),
	.aluifportOut_7(\ALU|aluif.portOut[7]~72_combout ),
	.dmemaddr6(\PR|dmemaddr~6_combout ),
	.aluifportOut_6(\ALU|aluif.portOut[6]~79_combout ),
	.dmemaddr7(\PR|dmemaddr~7_combout ),
	.aluifportOut_9(\ALU|aluif.portOut[9]~90_combout ),
	.dmemaddr8(\PR|dmemaddr~8_combout ),
	.aluifportOut_8(\ALU|aluif.portOut[8]~96_combout ),
	.dmemaddr9(\PR|dmemaddr~9_combout ),
	.aluifportOut_11(\ALU|aluif.portOut[11]~102_combout ),
	.dmemaddr10(\PR|dmemaddr~10_combout ),
	.aluifportOut_10(\ALU|aluif.portOut[10]~108_combout ),
	.dmemaddr11(\PR|dmemaddr~11_combout ),
	.aluifportOut_13(\ALU|aluif.portOut[13]~114_combout ),
	.dmemaddr12(\PR|dmemaddr~12_combout ),
	.aluifportOut_12(\ALU|aluif.portOut[12]~120_combout ),
	.dmemaddr13(\PR|dmemaddr~13_combout ),
	.aluifportOut_15(\ALU|aluif.portOut[15]~126_combout ),
	.dmemaddr14(\PR|dmemaddr~14_combout ),
	.aluifportOut_14(\ALU|aluif.portOut[14]~132_combout ),
	.dmemaddr15(\PR|dmemaddr~15_combout ),
	.aluifportOut_23(\ALU|aluif.portOut[23]~140_combout ),
	.dmemaddr16(\PR|dmemaddr~16_combout ),
	.aluifportOut_22(\ALU|aluif.portOut[22]~147_combout ),
	.dmemaddr17(\PR|dmemaddr~17_combout ),
	.aluifportOut_211(\ALU|aluif.portOut[21]~153_combout ),
	.dmemaddr18(\PR|dmemaddr~18_combout ),
	.aluifportOut_29(\ALU|aluif.portOut[29]~166_combout ),
	.dmemaddr19(\PR|dmemaddr~19_combout ),
	.prifpc_mem_29(\prif.pc_mem [29]),
	.aluifportOut_28(\ALU|aluif.portOut[28]~180_combout ),
	.dmemaddr20(\PR|dmemaddr~20_combout ),
	.prifpc_mem_28(\prif.pc_mem [28]),
	.aluifneg_flag(\ALU|aluif.neg_flag~19_combout ),
	.dmemaddr21(\PR|dmemaddr~21_combout ),
	.prifpc_mem_31(\prif.pc_mem [31]),
	.aluifportOut_30(\ALU|aluif.portOut[30]~189_combout ),
	.dmemaddr22(\PR|dmemaddr~22_combout ),
	.prifpc_mem_30(\prif.pc_mem [30]),
	.aluifportOut_20(\ALU|aluif.portOut[20]~195_combout ),
	.dmemaddr23(\PR|dmemaddr~23_combout ),
	.aluifportOut_17(\ALU|aluif.portOut[17]~201_combout ),
	.dmemaddr24(\PR|dmemaddr~24_combout ),
	.aluifportOut_16(\ALU|aluif.portOut[16]~207_combout ),
	.dmemaddr25(\PR|dmemaddr~25_combout ),
	.aluifportOut_19(\ALU|aluif.portOut[19]~213_combout ),
	.dmemaddr26(\PR|dmemaddr~26_combout ),
	.aluifportOut_18(\ALU|aluif.portOut[18]~221_combout ),
	.dmemaddr27(\PR|dmemaddr~27_combout ),
	.aluifportOut_25(\ALU|aluif.portOut[25]~234_combout ),
	.dmemaddr28(\PR|dmemaddr~28_combout ),
	.aluifportOut_24(\ALU|aluif.portOut[24]~241_combout ),
	.dmemaddr29(\PR|dmemaddr~29_combout ),
	.aluifportOut_27(\ALU|aluif.portOut[27]~249_combout ),
	.dmemaddr30(\PR|dmemaddr~30_combout ),
	.aluifportOut_26(\ALU|aluif.portOut[26]~257_combout ),
	.dmemaddr31(\PR|dmemaddr~31_combout ),
	.halt_mem(\PR|halt_mem~0_combout ),
	.dmemstore(\PR|dmemstore~0_combout ),
	.flush_idex(\HU|flush_idex~0_combout ),
	.Equal15(\CU|Equal15~0_combout ),
	.Equal11(\CU|Equal11~0_combout ),
	.Equal0(\CU|Equal0~0_combout ),
	.Equal10(\CU|Equal10~0_combout ),
	.Equal12(\CU|Equal12~0_combout ),
	.Equal20(\CU|Equal20~0_combout ),
	.Equal26(\CU|Equal26~0_combout ),
	.Equal25(\CU|Equal25~1_combout ),
	.Equal13(\CU|Equal13~0_combout ),
	.dataScr_ex(\PR|dataScr_ex~2_combout ),
	.WideNor0(\CU|WideNor0~2_combout ),
	.Selector0(\CU|Selector0~2_combout ),
	.ALUOP_ex(\PR|ALUOP_ex~0_combout ),
	.imm_ex(\PR|imm_ex~0_combout ),
	.ALUScr_ex(\PR|ALUScr_ex~11_combout ),
	.shamt_ex(\PR|shamt_ex~0_combout ),
	.ALUScr_ex1(\PR|ALUScr_ex~12_combout ),
	.Regwen_mem(\PR|Regwen_mem~0_combout ),
	.regwrite_mem(\PR|regwrite_mem~1_combout ),
	.regwrite_mem1(\PR|regwrite_mem~3_combout ),
	.regwrite_mem2(\PR|regwrite_mem~5_combout ),
	.regwrite_mem3(\PR|regwrite_mem~7_combout ),
	.regwrite_mem4(\PR|regwrite_mem~9_combout ),
	.rt_ex(\PR|rt_ex~0_combout ),
	.rt_ex1(\PR|rt_ex~1_combout ),
	.rt_ex2(\PR|rt_ex~2_combout ),
	.rt_ex3(\PR|rt_ex~3_combout ),
	.rt_ex4(\PR|rt_ex~4_combout ),
	.Regwen_wb(\PR|Regwen_wb~0_combout ),
	.regwrite_wb(\PR|regwrite_wb~0_combout ),
	.regwrite_wb1(\PR|regwrite_wb~1_combout ),
	.regwrite_wb2(\PR|regwrite_wb~2_combout ),
	.regwrite_wb3(\PR|regwrite_wb~3_combout ),
	.regwrite_wb4(\PR|regwrite_wb~4_combout ),
	.dmemload_wb(\PR|dmemload_wb~0_combout ),
	.dmemaddr_wb(\PR|dmemaddr_wb~0_combout ),
	.dataScr_wb(\PR|dataScr_wb~0_combout ),
	.dataScr_wb1(\PR|dataScr_wb~1_combout ),
	.prifpc_mem_1(\prif.pc_mem [1]),
	.pc_wb(\PR|pc_wb~0_combout ),
	.Mux622(\RF|Mux62~9_combout ),
	.Mux623(\RF|Mux62~19_combout ),
	.rdat2_ex(\PR|rdat2_ex~1_combout ),
	.prifrs_ex_01(\prif.rs_ex[0]~0_combout ),
	.prifrs_ex_11(\PR|prif.rs_ex[1]~0_combout ),
	.prifrs_ex_02(\PR|prif.rs_ex[0]~1_combout ),
	.prifrs_ex_31(\PR|prif.rs_ex[3]~2_combout ),
	.prifrs_ex_21(\PR|prif.rs_ex[2]~3_combout ),
	.prifrs_ex_41(\PR|prif.rs_ex[4]~4_combout ),
	.opcode_mem(\PR|opcode_mem~0_combout ),
	.opcode_mem1(\PR|opcode_mem~1_combout ),
	.opcode_mem2(\PR|opcode_mem~2_combout ),
	.opcode_mem3(\PR|opcode_mem~3_combout ),
	.opcode_mem4(\PR|opcode_mem~4_combout ),
	.opcode_mem5(\PR|opcode_mem~5_combout ),
	.Mux30(\RF|Mux30~9_combout ),
	.Mux301(\RF|Mux30~19_combout ),
	.rdat1_ex(\PR|rdat1_ex~1_combout ),
	.imm_ex1(\PR|imm_ex~1_combout ),
	.shamt_ex1(\PR|shamt_ex~1_combout ),
	.dmemload_wb1(\PR|dmemload_wb~1_combout ),
	.dmemaddr_wb1(\PR|dmemaddr_wb~1_combout ),
	.prifpc_mem_0(\prif.pc_mem [0]),
	.pc_wb1(\PR|pc_wb~1_combout ),
	.Mux632(\RF|Mux63~9_combout ),
	.Mux633(\RF|Mux63~19_combout ),
	.rdat2_ex1(\PR|rdat2_ex~3_combout ),
	.Mux31(\RF|Mux31~9_combout ),
	.Mux311(\RF|Mux31~19_combout ),
	.rdat1_ex1(\PR|rdat1_ex~3_combout ),
	.dmemload_wb2(\PR|dmemload_wb~2_combout ),
	.dmemaddr_wb2(\PR|dmemaddr_wb~2_combout ),
	.prifpc_mem_3(\prif.pc_mem [3]),
	.pc_wb2(\PR|pc_wb~2_combout ),
	.Mux60(\RF|Mux60~9_combout ),
	.Mux601(\RF|Mux60~19_combout ),
	.rdat2_ex2(\PR|rdat2_ex~5_combout ),
	.imm_ex2(\PR|imm_ex~2_combout ),
	.shamt_ex2(\PR|shamt_ex~2_combout ),
	.imm_ex3(\PR|imm_ex~3_combout ),
	.shamt_ex3(\PR|shamt_ex~3_combout ),
	.dmemload_wb3(\PR|dmemload_wb~3_combout ),
	.dmemaddr_wb3(\PR|dmemaddr_wb~3_combout ),
	.prifpc_mem_2(\prif.pc_mem [2]),
	.pc_wb3(\PR|pc_wb~3_combout ),
	.Mux611(\RF|Mux61~9_combout ),
	.Mux612(\RF|Mux61~19_combout ),
	.rdat2_ex3(\PR|rdat2_ex~7_combout ),
	.dmemload_wb4(\PR|dmemload_wb~4_combout ),
	.dmemaddr_wb4(\PR|dmemaddr_wb~4_combout ),
	.prifpc_mem_4(\prif.pc_mem [4]),
	.pc_wb4(\PR|pc_wb~4_combout ),
	.Mux59(\RF|Mux59~9_combout ),
	.Mux591(\RF|Mux59~19_combout ),
	.rdat2_ex4(\PR|rdat2_ex~9_combout ),
	.imm_ex4(\PR|imm_ex~4_combout ),
	.shamt_ex4(\PR|shamt_ex~4_combout ),
	.instr_ex(\PR|instr_ex~0_combout ),
	.dmemload_wb5(\PR|dmemload_wb~5_combout ),
	.imm_wb(\PR|imm_wb~0_combout ),
	.dmemaddr_wb5(\PR|dmemaddr_wb~5_combout ),
	.pc_wb5(\PR|pc_wb~5_combout ),
	.Mux321(\RF|Mux32~9_combout ),
	.Mux322(\RF|Mux32~19_combout ),
	.rdat2_ex5(\PR|rdat2_ex~11_combout ),
	.imm_mem(\PR|imm_mem~0_combout ),
	.imm_wb1(\PR|imm_wb~1_combout ),
	.dmemload_wb6(\PR|dmemload_wb~6_combout ),
	.dmemaddr_wb6(\PR|dmemaddr_wb~6_combout ),
	.pc_wb6(\PR|pc_wb~6_combout ),
	.Mux331(\RF|Mux33~9_combout ),
	.Mux332(\RF|Mux33~19_combout ),
	.rdat2_ex6(\PR|rdat2_ex~13_combout ),
	.imm_mem1(\PR|imm_mem~1_combout ),
	.dmemload_wb7(\PR|dmemload_wb~7_combout ),
	.imm_wb2(\PR|imm_wb~2_combout ),
	.dmemaddr_wb7(\PR|dmemaddr_wb~7_combout ),
	.pc_wb7(\PR|pc_wb~7_combout ),
	.Mux341(\RF|Mux34~9_combout ),
	.Mux342(\RF|Mux34~19_combout ),
	.rdat2_ex7(\PR|rdat2_ex~15_combout ),
	.imm_mem2(\PR|imm_mem~2_combout ),
	.imm_ex5(\PR|imm_ex~5_combout ),
	.dmemload_wb8(\PR|dmemload_wb~8_combout ),
	.dmemaddr_wb8(\PR|dmemaddr_wb~8_combout ),
	.prifpc_mem_5(\prif.pc_mem [5]),
	.pc_wb8(\PR|pc_wb~8_combout ),
	.Mux58(\RF|Mux58~9_combout ),
	.Mux581(\RF|Mux58~19_combout ),
	.rdat2_ex8(\PR|rdat2_ex~17_combout ),
	.imm_ex6(\PR|imm_ex~6_combout ),
	.dmemload_wb9(\PR|dmemload_wb~9_combout ),
	.dmemaddr_wb9(\PR|dmemaddr_wb~9_combout ),
	.prifpc_mem_15(\prif.pc_mem [15]),
	.pc_wb9(\PR|pc_wb~9_combout ),
	.Mux48(\RF|Mux48~9_combout ),
	.Mux481(\RF|Mux48~19_combout ),
	.rdat2_ex9(\PR|rdat2_ex~19_combout ),
	.imm_ex7(\PR|imm_ex~7_combout ),
	.dmemload_wb10(\PR|dmemload_wb~10_combout ),
	.dmemaddr_wb10(\PR|dmemaddr_wb~10_combout ),
	.prifpc_mem_14(\prif.pc_mem [14]),
	.pc_wb10(\PR|pc_wb~10_combout ),
	.Mux49(\RF|Mux49~9_combout ),
	.Mux491(\RF|Mux49~19_combout ),
	.rdat2_ex10(\PR|rdat2_ex~21_combout ),
	.imm_ex8(\PR|imm_ex~8_combout ),
	.dmemload_wb11(\PR|dmemload_wb~11_combout ),
	.dmemaddr_wb11(\PR|dmemaddr_wb~11_combout ),
	.prifpc_mem_13(\prif.pc_mem [13]),
	.pc_wb11(\PR|pc_wb~11_combout ),
	.Mux50(\RF|Mux50~9_combout ),
	.Mux501(\RF|Mux50~19_combout ),
	.rdat2_ex11(\PR|rdat2_ex~23_combout ),
	.imm_ex9(\PR|imm_ex~9_combout ),
	.dmemload_wb12(\PR|dmemload_wb~12_combout ),
	.dmemaddr_wb12(\PR|dmemaddr_wb~12_combout ),
	.prifpc_mem_12(\prif.pc_mem [12]),
	.pc_wb12(\PR|pc_wb~12_combout ),
	.Mux51(\RF|Mux51~9_combout ),
	.Mux511(\RF|Mux51~19_combout ),
	.rdat2_ex12(\PR|rdat2_ex~25_combout ),
	.imm_ex10(\PR|imm_ex~10_combout ),
	.dmemload_wb13(\PR|dmemload_wb~13_combout ),
	.dmemaddr_wb13(\PR|dmemaddr_wb~13_combout ),
	.prifpc_mem_11(\prif.pc_mem [11]),
	.pc_wb13(\PR|pc_wb~13_combout ),
	.Mux52(\RF|Mux52~9_combout ),
	.Mux521(\RF|Mux52~19_combout ),
	.rdat2_ex13(\PR|rdat2_ex~27_combout ),
	.imm_ex11(\PR|imm_ex~11_combout ),
	.dmemload_wb14(\PR|dmemload_wb~14_combout ),
	.dmemaddr_wb14(\PR|dmemaddr_wb~14_combout ),
	.prifpc_mem_10(\prif.pc_mem [10]),
	.pc_wb14(\PR|pc_wb~14_combout ),
	.Mux53(\RF|Mux53~9_combout ),
	.Mux531(\RF|Mux53~19_combout ),
	.rdat2_ex14(\PR|rdat2_ex~29_combout ),
	.imm_ex12(\PR|imm_ex~12_combout ),
	.dmemload_wb15(\PR|dmemload_wb~15_combout ),
	.dmemaddr_wb15(\PR|dmemaddr_wb~15_combout ),
	.prifpc_mem_9(\prif.pc_mem [9]),
	.pc_wb15(\PR|pc_wb~15_combout ),
	.Mux54(\RF|Mux54~9_combout ),
	.Mux541(\RF|Mux54~19_combout ),
	.rdat2_ex15(\PR|rdat2_ex~31_combout ),
	.imm_ex13(\PR|imm_ex~13_combout ),
	.dmemload_wb16(\PR|dmemload_wb~16_combout ),
	.dmemaddr_wb16(\PR|dmemaddr_wb~16_combout ),
	.prifpc_mem_6(\prif.pc_mem [6]),
	.pc_wb16(\PR|pc_wb~16_combout ),
	.Mux57(\RF|Mux57~9_combout ),
	.Mux571(\RF|Mux57~19_combout ),
	.rdat2_ex16(\PR|rdat2_ex~33_combout ),
	.dmemload_wb17(\PR|dmemload_wb~17_combout ),
	.imm_wb3(\PR|imm_wb~3_combout ),
	.dmemaddr_wb17(\PR|dmemaddr_wb~17_combout ),
	.prifpc_mem_27(\prif.pc_mem [27]),
	.pc_wb17(\PR|pc_wb~17_combout ),
	.Mux361(\RF|Mux36~9_combout ),
	.Mux362(\RF|Mux36~19_combout ),
	.rdat2_ex17(\PR|rdat2_ex~35_combout ),
	.imm_mem3(\PR|imm_mem~3_combout ),
	.dmemload_wb18(\PR|dmemload_wb~18_combout ),
	.imm_wb4(\PR|imm_wb~4_combout ),
	.dmemaddr_wb18(\PR|dmemaddr_wb~18_combout ),
	.prifpc_mem_23(\prif.pc_mem [23]),
	.pc_wb18(\PR|pc_wb~18_combout ),
	.Mux401(\RF|Mux40~9_combout ),
	.Mux402(\RF|Mux40~19_combout ),
	.rdat2_ex18(\PR|rdat2_ex~37_combout ),
	.imm_mem4(\PR|imm_mem~4_combout ),
	.imm_wb5(\PR|imm_wb~5_combout ),
	.dmemload_wb19(\PR|dmemload_wb~19_combout ),
	.dmemaddr_wb19(\PR|dmemaddr_wb~19_combout ),
	.prifpc_mem_18(\prif.pc_mem [18]),
	.pc_wb19(\PR|pc_wb~19_combout ),
	.Mux451(\RF|Mux45~9_combout ),
	.Mux452(\RF|Mux45~19_combout ),
	.rdat2_ex19(\PR|rdat2_ex~39_combout ),
	.imm_mem5(\PR|imm_mem~5_combout ),
	.imm_wb6(\PR|imm_wb~6_combout ),
	.dmemload_wb20(\PR|dmemload_wb~20_combout ),
	.dmemaddr_wb20(\PR|dmemaddr_wb~20_combout ),
	.prifpc_mem_24(\prif.pc_mem [24]),
	.pc_wb20(\PR|pc_wb~20_combout ),
	.Mux391(\RF|Mux39~9_combout ),
	.Mux392(\RF|Mux39~19_combout ),
	.rdat2_ex20(\PR|rdat2_ex~41_combout ),
	.imm_mem6(\PR|imm_mem~6_combout ),
	.imm_wb7(\PR|imm_wb~7_combout ),
	.dmemload_wb21(\PR|dmemload_wb~21_combout ),
	.dmemaddr_wb21(\PR|dmemaddr_wb~21_combout ),
	.prifpc_mem_16(\prif.pc_mem [16]),
	.pc_wb21(\PR|pc_wb~21_combout ),
	.Mux471(\RF|Mux47~9_combout ),
	.Mux472(\RF|Mux47~19_combout ),
	.rdat2_ex21(\PR|rdat2_ex~43_combout ),
	.imm_mem7(\PR|imm_mem~7_combout ),
	.dmemload_wb22(\PR|dmemload_wb~22_combout ),
	.imm_wb8(\PR|imm_wb~8_combout ),
	.dmemaddr_wb22(\PR|dmemaddr_wb~22_combout ),
	.prifpc_mem_19(\prif.pc_mem [19]),
	.pc_wb22(\PR|pc_wb~22_combout ),
	.Mux441(\RF|Mux44~9_combout ),
	.Mux442(\RF|Mux44~19_combout ),
	.rdat2_ex22(\PR|rdat2_ex~45_combout ),
	.imm_mem8(\PR|imm_mem~8_combout ),
	.dmemload_wb23(\PR|dmemload_wb~23_combout ),
	.imm_wb9(\PR|imm_wb~9_combout ),
	.dmemaddr_wb23(\PR|dmemaddr_wb~23_combout ),
	.prifpc_mem_17(\prif.pc_mem [17]),
	.pc_wb23(\PR|pc_wb~23_combout ),
	.Mux461(\RF|Mux46~9_combout ),
	.Mux462(\RF|Mux46~19_combout ),
	.rdat2_ex23(\PR|rdat2_ex~47_combout ),
	.imm_mem9(\PR|imm_mem~9_combout ),
	.dmemload_wb24(\PR|dmemload_wb~24_combout ),
	.imm_wb10(\PR|imm_wb~10_combout ),
	.dmemaddr_wb24(\PR|dmemaddr_wb~24_combout ),
	.prifpc_mem_21(\prif.pc_mem [21]),
	.pc_wb24(\PR|pc_wb~24_combout ),
	.Mux421(\RF|Mux42~9_combout ),
	.Mux422(\RF|Mux42~19_combout ),
	.rdat2_ex24(\PR|rdat2_ex~49_combout ),
	.imm_mem10(\PR|imm_mem~10_combout ),
	.imm_wb11(\PR|imm_wb~11_combout ),
	.dmemload_wb25(\PR|dmemload_wb~25_combout ),
	.dmemaddr_wb25(\PR|dmemaddr_wb~25_combout ),
	.prifpc_mem_20(\prif.pc_mem [20]),
	.pc_wb25(\PR|pc_wb~25_combout ),
	.Mux431(\RF|Mux43~9_combout ),
	.Mux432(\RF|Mux43~19_combout ),
	.rdat2_ex25(\PR|rdat2_ex~51_combout ),
	.imm_mem11(\PR|imm_mem~11_combout ),
	.imm_wb12(\PR|imm_wb~12_combout ),
	.dmemload_wb26(\PR|dmemload_wb~26_combout ),
	.dmemaddr_wb26(\PR|dmemaddr_wb~26_combout ),
	.pc_wb26(\PR|pc_wb~26_combout ),
	.Mux351(\RF|Mux35~9_combout ),
	.Mux352(\RF|Mux35~19_combout ),
	.rdat2_ex26(\PR|rdat2_ex~53_combout ),
	.imm_mem12(\PR|imm_mem~12_combout ),
	.imm_wb13(\PR|imm_wb~13_combout ),
	.dmemload_wb27(\PR|dmemload_wb~27_combout ),
	.dmemaddr_wb27(\PR|dmemaddr_wb~27_combout ),
	.prifpc_mem_26(\prif.pc_mem [26]),
	.pc_wb27(\PR|pc_wb~27_combout ),
	.Mux371(\RF|Mux37~9_combout ),
	.Mux372(\RF|Mux37~19_combout ),
	.rdat2_ex27(\PR|rdat2_ex~55_combout ),
	.imm_mem13(\PR|imm_mem~13_combout ),
	.imm_ex14(\PR|imm_ex~14_combout ),
	.dmemload_wb28(\PR|dmemload_wb~28_combout ),
	.dmemaddr_wb28(\PR|dmemaddr_wb~28_combout ),
	.prifpc_mem_8(\prif.pc_mem [8]),
	.pc_wb28(\PR|pc_wb~28_combout ),
	.Mux55(\RF|Mux55~9_combout ),
	.Mux551(\RF|Mux55~19_combout ),
	.rdat2_ex28(\PR|rdat2_ex~57_combout ),
	.imm_ex15(\PR|imm_ex~15_combout ),
	.dmemload_wb29(\PR|dmemload_wb~29_combout ),
	.dmemaddr_wb29(\PR|dmemaddr_wb~29_combout ),
	.prifpc_mem_7(\prif.pc_mem [7]),
	.pc_wb29(\PR|pc_wb~29_combout ),
	.Mux56(\RF|Mux56~9_combout ),
	.Mux561(\RF|Mux56~19_combout ),
	.rdat2_ex29(\PR|rdat2_ex~59_combout ),
	.imm_wb14(\PR|imm_wb~14_combout ),
	.dmemload_wb30(\PR|dmemload_wb~30_combout ),
	.dmemaddr_wb30(\PR|dmemaddr_wb~30_combout ),
	.prifpc_mem_22(\prif.pc_mem [22]),
	.pc_wb30(\PR|pc_wb~30_combout ),
	.Mux411(\RF|Mux41~9_combout ),
	.Mux412(\RF|Mux41~19_combout ),
	.rdat2_ex30(\PR|rdat2_ex~61_combout ),
	.imm_mem14(\PR|imm_mem~14_combout ),
	.dmemload_wb31(\PR|dmemload_wb~31_combout ),
	.imm_wb15(\PR|imm_wb~15_combout ),
	.dmemaddr_wb31(\PR|dmemaddr_wb~31_combout ),
	.prifpc_mem_25(\prif.pc_mem [25]),
	.pc_wb31(\PR|pc_wb~31_combout ),
	.Mux381(\RF|Mux38~9_combout ),
	.Mux382(\RF|Mux38~19_combout ),
	.rdat2_ex31(\PR|rdat2_ex~63_combout ),
	.imm_mem15(\PR|imm_mem~15_combout ),
	.Equal4(\CU|Equal4~0_combout ),
	.ALUOP_ex1(\PR|ALUOP_ex~2_combout ),
	.Selector2(\CU|Selector2~4_combout ),
	.Selector21(\CU|Selector2~5_combout ),
	.ALUOP_ex2(\PR|ALUOP_ex~3_combout ),
	.Mux29(\RF|Mux29~9_combout ),
	.Mux291(\RF|Mux29~19_combout ),
	.rdat1_ex2(\PR|rdat1_ex~5_combout ),
	.Mux27(\RF|Mux27~9_combout ),
	.Mux271(\RF|Mux27~19_combout ),
	.rdat1_ex3(\PR|rdat1_ex~7_combout ),
	.Mux28(\RF|Mux28~9_combout ),
	.Mux281(\RF|Mux28~19_combout ),
	.rdat1_ex4(\PR|rdat1_ex~9_combout ),
	.Mux23(\RF|Mux23~9_combout ),
	.Mux231(\RF|Mux23~19_combout ),
	.rdat1_ex5(\PR|rdat1_ex~11_combout ),
	.Mux24(\RF|Mux24~9_combout ),
	.Mux241(\RF|Mux24~19_combout ),
	.rdat1_ex6(\PR|rdat1_ex~13_combout ),
	.Mux25(\RF|Mux25~9_combout ),
	.Mux251(\RF|Mux25~19_combout ),
	.rdat1_ex7(\PR|rdat1_ex~15_combout ),
	.Mux26(\RF|Mux26~9_combout ),
	.Mux261(\RF|Mux26~19_combout ),
	.rdat1_ex8(\PR|rdat1_ex~17_combout ),
	.Mux15(\RF|Mux15~9_combout ),
	.Mux151(\RF|Mux15~19_combout ),
	.rdat1_ex9(\PR|rdat1_ex~19_combout ),
	.Mux16(\RF|Mux16~9_combout ),
	.Mux161(\RF|Mux16~19_combout ),
	.rdat1_ex10(\PR|rdat1_ex~21_combout ),
	.Mux17(\RF|Mux17~9_combout ),
	.Mux171(\RF|Mux17~19_combout ),
	.rdat1_ex11(\PR|rdat1_ex~23_combout ),
	.Mux18(\RF|Mux18~9_combout ),
	.Mux181(\RF|Mux18~19_combout ),
	.rdat1_ex12(\PR|rdat1_ex~25_combout ),
	.Mux20(\RF|Mux20~9_combout ),
	.Mux201(\RF|Mux20~19_combout ),
	.rdat1_ex13(\PR|rdat1_ex~27_combout ),
	.Mux19(\RF|Mux19~9_combout ),
	.Mux191(\RF|Mux19~19_combout ),
	.rdat1_ex14(\PR|rdat1_ex~29_combout ),
	.Mux21(\RF|Mux21~9_combout ),
	.Mux211(\RF|Mux21~19_combout ),
	.rdat1_ex15(\PR|rdat1_ex~31_combout ),
	.Mux22(\RF|Mux22~9_combout ),
	.Mux221(\RF|Mux22~19_combout ),
	.rdat1_ex16(\PR|rdat1_ex~33_combout ),
	.Mux13(\RF|Mux13~9_combout ),
	.Mux131(\RF|Mux13~19_combout ),
	.rdat1_ex17(\PR|rdat1_ex~35_combout ),
	.Mux14(\RF|Mux14~9_combout ),
	.Mux141(\RF|Mux14~19_combout ),
	.rdat1_ex18(\PR|rdat1_ex~37_combout ),
	.Mux11(\RF|Mux11~9_combout ),
	.Mux111(\RF|Mux11~19_combout ),
	.rdat1_ex19(\PR|rdat1_ex~39_combout ),
	.Mux12(\RF|Mux12~9_combout ),
	.Mux121(\RF|Mux12~19_combout ),
	.rdat1_ex20(\PR|rdat1_ex~41_combout ),
	.Mux9(\RF|Mux9~9_combout ),
	.Mux91(\RF|Mux9~19_combout ),
	.rdat1_ex21(\PR|rdat1_ex~43_combout ),
	.Mux10(\RF|Mux10~9_combout ),
	.Mux101(\RF|Mux10~19_combout ),
	.rdat1_ex22(\PR|rdat1_ex~45_combout ),
	.Mux7(\RF|Mux7~9_combout ),
	.Mux71(\RF|Mux7~19_combout ),
	.rdat1_ex23(\PR|rdat1_ex~47_combout ),
	.Mux8(\RF|Mux8~9_combout ),
	.Mux81(\RF|Mux8~19_combout ),
	.rdat1_ex24(\PR|rdat1_ex~49_combout ),
	.Mux0(\RF|Mux0~9_combout ),
	.Mux01(\RF|Mux0~19_combout ),
	.rdat1_ex25(\PR|rdat1_ex~51_combout ),
	.Mux1(\RF|Mux1~9_combout ),
	.Mux110(\RF|Mux1~19_combout ),
	.rdat1_ex26(\PR|rdat1_ex~53_combout ),
	.Mux2(\RF|Mux2~9_combout ),
	.Mux210(\RF|Mux2~19_combout ),
	.rdat1_ex27(\PR|rdat1_ex~55_combout ),
	.Mux5(\RF|Mux5~9_combout ),
	.Mux510(\RF|Mux5~19_combout ),
	.rdat1_ex28(\PR|rdat1_ex~57_combout ),
	.Mux6(\RF|Mux6~9_combout ),
	.Mux64(\RF|Mux6~19_combout ),
	.rdat1_ex29(\PR|rdat1_ex~59_combout ),
	.Mux3(\RF|Mux3~9_combout ),
	.Mux310(\RF|Mux3~19_combout ),
	.rdat1_ex30(\PR|rdat1_ex~61_combout ),
	.Mux4(\RF|Mux4~9_combout ),
	.Mux410(\RF|Mux4~19_combout ),
	.rdat1_ex31(\PR|rdat1_ex~63_combout ),
	.ALUScr_ex2(\PR|ALUScr_ex~13_combout ),
	.Selector3(\CU|Selector3~5_combout ),
	.ALUOP_ex3(\PR|ALUOP_ex~4_combout ),
	.aluifportOut_53(\ALU|aluif.portOut[5]~258_combout ),
	.instr_mem(\PR|instr_mem~0_combout ),
	.instr_mem1(\PR|instr_mem~1_combout ),
	.instr_mem2(\PR|instr_mem~2_combout ),
	.instr_mem3(\PR|instr_mem~3_combout ),
	.instr_mem4(\PR|instr_mem~4_combout ),
	.instr_mem5(\PR|instr_mem~5_combout ),
	.rdat1_mem(\PR|rdat1_mem~0_combout ),
	.PCScr_mem(\PR|PCScr_mem~0_combout ),
	.pc_bran_mem(\PR|pc_bran_mem~0_combout ),
	.PCScr_mem1(\PR|PCScr_mem~1_combout ),
	.opcode_ex(\PR|opcode_ex~0_combout ),
	.opcode_ex1(\PR|opcode_ex~1_combout ),
	.opcode_ex2(\PR|opcode_ex~2_combout ),
	.opcode_ex3(\PR|opcode_ex~3_combout ),
	.opcode_ex4(\PR|opcode_ex~4_combout ),
	.Equal131(\CU|Equal13~1_combout ),
	.memren_ex(\PR|memren_ex~0_combout ),
	.memwen_ex(\PR|memwen_ex~0_combout ),
	.rdat1_mem1(\PR|rdat1_mem~1_combout ),
	.pc_bran_mem1(\PR|pc_bran_mem~1_combout ),
	.rdat1_mem2(\PR|rdat1_mem~2_combout ),
	.pc_bran_mem2(\PR|pc_bran_mem~2_combout ),
	.rdat1_mem3(\PR|rdat1_mem~3_combout ),
	.pc_bran_mem3(\PR|pc_bran_mem~3_combout ),
	.rdat1_mem4(\PR|rdat1_mem~4_combout ),
	.pc_bran_mem4(\PR|pc_bran_mem~4_combout ),
	.rdat1_mem5(\PR|rdat1_mem~5_combout ),
	.pc_bran_mem5(\PR|pc_bran_mem~5_combout ),
	.rdat1_mem6(\PR|rdat1_mem~6_combout ),
	.pc_bran_mem6(\PR|pc_bran_mem~6_combout ),
	.rdat1_mem7(\PR|rdat1_mem~7_combout ),
	.pc_bran_mem7(\PR|pc_bran_mem~7_combout ),
	.rdat1_mem8(\PR|rdat1_mem~8_combout ),
	.pc_bran_mem8(\PR|pc_bran_mem~8_combout ),
	.instr_mem6(\PR|instr_mem~6_combout ),
	.rdat1_mem9(\PR|rdat1_mem~9_combout ),
	.pc_bran_mem9(\PR|pc_bran_mem~9_combout ),
	.instr_mem7(\PR|instr_mem~7_combout ),
	.rdat1_mem10(\PR|rdat1_mem~10_combout ),
	.pc_bran_mem10(\PR|pc_bran_mem~10_combout ),
	.instr_mem8(\PR|instr_mem~8_combout ),
	.rdat1_mem11(\PR|rdat1_mem~11_combout ),
	.pc_bran_mem11(\PR|pc_bran_mem~11_combout ),
	.instr_mem9(\PR|instr_mem~9_combout ),
	.rdat1_mem12(\PR|rdat1_mem~12_combout ),
	.pc_bran_mem12(\PR|pc_bran_mem~12_combout ),
	.instr_mem10(\PR|instr_mem~10_combout ),
	.rdat1_mem13(\PR|rdat1_mem~13_combout ),
	.pc_bran_mem13(\PR|pc_bran_mem~13_combout ),
	.instr_mem11(\PR|instr_mem~11_combout ),
	.rdat1_mem14(\PR|rdat1_mem~14_combout ),
	.pc_bran_mem14(\PR|pc_bran_mem~14_combout ),
	.instr_mem12(\PR|instr_mem~12_combout ),
	.rdat1_mem15(\PR|rdat1_mem~15_combout ),
	.pc_bran_mem15(\PR|pc_bran_mem~15_combout ),
	.instr_mem13(\PR|instr_mem~13_combout ),
	.rdat1_mem16(\PR|rdat1_mem~16_combout ),
	.pc_bran_mem16(\PR|pc_bran_mem~16_combout ),
	.instr_mem14(\PR|instr_mem~14_combout ),
	.rdat1_mem17(\PR|rdat1_mem~17_combout ),
	.pc_bran_mem17(\PR|pc_bran_mem~17_combout ),
	.instr_mem15(\PR|instr_mem~15_combout ),
	.rdat1_mem18(\PR|rdat1_mem~18_combout ),
	.pc_bran_mem18(\PR|pc_bran_mem~18_combout ),
	.instr_mem16(\PR|instr_mem~16_combout ),
	.rdat1_mem19(\PR|rdat1_mem~19_combout ),
	.pc_bran_mem19(\PR|pc_bran_mem~19_combout ),
	.prifpc_mem_151(\prif.pc_mem[15]~0_combout ),
	.prifpc_mem_291(\PR|prif.pc_mem[29]~0_combout ),
	.rdat1_mem20(\PR|rdat1_mem~20_combout ),
	.pc_bran_mem20(\PR|pc_bran_mem~20_combout ),
	.prifpc_mem_281(\PR|prif.pc_mem[28]~1_combout ),
	.rdat1_mem21(\PR|rdat1_mem~21_combout ),
	.pc_bran_mem21(\PR|pc_bran_mem~21_combout ),
	.prifpc_mem_311(\PR|prif.pc_mem[31]~2_combout ),
	.rdat1_mem22(\PR|rdat1_mem~22_combout ),
	.pc_bran_mem22(\PR|pc_bran_mem~22_combout ),
	.prifpc_mem_301(\PR|prif.pc_mem[30]~3_combout ),
	.rdat1_mem23(\PR|rdat1_mem~23_combout ),
	.pc_bran_mem23(\PR|pc_bran_mem~23_combout ),
	.instr_mem17(\PR|instr_mem~17_combout ),
	.rdat1_mem24(\PR|rdat1_mem~24_combout ),
	.pc_bran_mem24(\PR|pc_bran_mem~24_combout ),
	.instr_mem18(\PR|instr_mem~18_combout ),
	.rdat1_mem25(\PR|rdat1_mem~25_combout ),
	.pc_bran_mem25(\PR|pc_bran_mem~25_combout ),
	.instr_mem19(\PR|instr_mem~19_combout ),
	.rdat1_mem26(\PR|rdat1_mem~26_combout ),
	.pc_bran_mem26(\PR|pc_bran_mem~26_combout ),
	.instr_mem20(\PR|instr_mem~20_combout ),
	.rdat1_mem27(\PR|rdat1_mem~27_combout ),
	.pc_bran_mem27(\PR|pc_bran_mem~27_combout ),
	.instr_mem21(\PR|instr_mem~21_combout ),
	.rdat1_mem28(\PR|rdat1_mem~28_combout ),
	.pc_bran_mem28(\PR|pc_bran_mem~28_combout ),
	.instr_mem22(\PR|instr_mem~22_combout ),
	.rdat1_mem29(\PR|rdat1_mem~29_combout ),
	.pc_bran_mem29(\PR|pc_bran_mem~29_combout ),
	.instr_mem23(\PR|instr_mem~23_combout ),
	.rdat1_mem30(\PR|rdat1_mem~30_combout ),
	.pc_bran_mem30(\PR|pc_bran_mem~30_combout ),
	.instr_mem24(\PR|instr_mem~24_combout ),
	.rdat1_mem31(\PR|rdat1_mem~31_combout ),
	.pc_bran_mem31(\PR|pc_bran_mem~31_combout ),
	.instr_mem25(\PR|instr_mem~25_combout ),
	.dmemstore1(\PR|dmemstore~1_combout ),
	.dmemstore2(\PR|dmemstore~2_combout ),
	.Mux602(\Mux60~1_combout ),
	.dmemstore3(\PR|dmemstore~3_combout ),
	.Mux592(\Mux59~1_combout ),
	.dmemstore4(\PR|dmemstore~4_combout ),
	.Mux582(\Mux58~1_combout ),
	.dmemstore5(\PR|dmemstore~5_combout ),
	.Mux572(\Mux57~1_combout ),
	.dmemstore6(\PR|dmemstore~6_combout ),
	.Mux562(\Mux56~1_combout ),
	.dmemstore7(\PR|dmemstore~7_combout ),
	.Mux552(\Mux55~1_combout ),
	.dmemstore8(\PR|dmemstore~8_combout ),
	.Mux542(\Mux54~1_combout ),
	.dmemstore9(\PR|dmemstore~9_combout ),
	.Mux532(\Mux53~1_combout ),
	.dmemstore10(\PR|dmemstore~10_combout ),
	.Mux522(\Mux52~1_combout ),
	.dmemstore11(\PR|dmemstore~11_combout ),
	.Mux512(\Mux51~1_combout ),
	.dmemstore12(\PR|dmemstore~12_combout ),
	.Mux502(\Mux50~1_combout ),
	.dmemstore13(\PR|dmemstore~13_combout ),
	.Mux492(\Mux49~1_combout ),
	.dmemstore14(\PR|dmemstore~14_combout ),
	.Mux482(\Mux48~1_combout ),
	.dmemstore15(\PR|dmemstore~15_combout ),
	.dmemstore16(\PR|dmemstore~16_combout ),
	.dmemstore17(\PR|dmemstore~17_combout ),
	.dmemstore18(\PR|dmemstore~18_combout ),
	.dmemstore19(\PR|dmemstore~19_combout ),
	.dmemstore20(\PR|dmemstore~20_combout ),
	.dmemstore21(\PR|dmemstore~21_combout ),
	.dmemstore22(\PR|dmemstore~22_combout ),
	.dmemstore23(\PR|dmemstore~23_combout ),
	.dmemstore24(\PR|dmemstore~24_combout ),
	.dmemstore25(\PR|dmemstore~25_combout ),
	.dmemstore26(\PR|dmemstore~26_combout ),
	.dmemstore27(\PR|dmemstore~27_combout ),
	.dmemstore28(\PR|dmemstore~28_combout ),
	.dmemstore29(\PR|dmemstore~29_combout ),
	.dmemstore30(\PR|dmemstore~30_combout ),
	.dmemstore31(\PR|dmemstore~31_combout ),
	.halt_ex(\PR|halt_ex~0_combout ),
	.prifhalt_wb(\prif.halt_wb~q ),
	.ifid_en(\HU|ifid_en~1_combout ),
	.imemload_id(\PR|imemload_id~0_combout ),
	.imemload_id1(\PR|imemload_id~1_combout ),
	.imemload_id2(\PR|imemload_id~2_combout ),
	.imemload_id3(\PR|imemload_id~3_combout ),
	.imemload_id4(\PR|imemload_id~4_combout ),
	.imemload_id5(\PR|imemload_id~5_combout ),
	.imemload_id6(\PR|imemload_id~6_combout ),
	.imemload_id7(\PR|imemload_id~7_combout ),
	.imemload_id8(\PR|imemload_id~8_combout ),
	.imemload_id9(\PR|imemload_id~9_combout ),
	.imemload_id10(\PR|imemload_id~10_combout ),
	.imemload_id11(\PR|imemload_id~11_combout ),
	.imemload_id12(\PR|imemload_id~12_combout ),
	.Regwen_ex(\PR|Regwen_ex~0_combout ),
	.rd_ex(\PR|rd_ex~0_combout ),
	.RegDest_ex(\PR|RegDest_ex~0_combout ),
	.RegDest_ex1(\PR|RegDest_ex~1_combout ),
	.rd_ex1(\PR|rd_ex~1_combout ),
	.rd_ex2(\PR|rd_ex~2_combout ),
	.rd_ex3(\PR|rd_ex~3_combout ),
	.rd_ex4(\PR|rd_ex~4_combout ),
	.imemload_id13(\PR|imemload_id~13_combout ),
	.imemload_id14(\PR|imemload_id~14_combout ),
	.imemload_id15(\PR|imemload_id~15_combout ),
	.imemload_id16(\PR|imemload_id~16_combout ),
	.imemload_id17(\PR|imemload_id~17_combout ),
	.dataScr_mem(\PR|dataScr_mem~0_combout ),
	.dataScr_mem1(\PR|dataScr_mem~1_combout ),
	.prifpc_mem_110(\PR|prif.pc_mem[1]~4_combout ),
	.imemload_id18(\PR|imemload_id~18_combout ),
	.imemload_id19(\PR|imemload_id~19_combout ),
	.imemload_id20(\PR|imemload_id~20_combout ),
	.imemload_id21(\PR|imemload_id~21_combout ),
	.imemload_id22(\PR|imemload_id~22_combout ),
	.opcode_ex5(\PR|opcode_ex~5_combout ),
	.imemload_id23(\PR|imemload_id~23_combout ),
	.prifpc_mem_01(\PR|prif.pc_mem[0]~5_combout ),
	.prifpc_mem_32(\PR|prif.pc_mem[3]~6_combout ),
	.imemload_id24(\PR|imemload_id~24_combout ),
	.imemload_id25(\PR|imemload_id~25_combout ),
	.prifpc_mem_210(\PR|prif.pc_mem[2]~7_combout ),
	.prifpc_mem_41(\PR|prif.pc_mem[4]~8_combout ),
	.imemload_id26(\PR|imemload_id~26_combout ),
	.imemload_id27(\PR|imemload_id~27_combout ),
	.prifpc_mem_51(\PR|prif.pc_mem[5]~9_combout ),
	.prifpc_mem_152(\PR|prif.pc_mem[15]~10_combout ),
	.imemload_id28(\PR|imemload_id~28_combout ),
	.prifpc_mem_141(\PR|prif.pc_mem[14]~11_combout ),
	.imemload_id29(\PR|imemload_id~29_combout ),
	.prifpc_mem_131(\PR|prif.pc_mem[13]~12_combout ),
	.imemload_id30(\PR|imemload_id~30_combout ),
	.prifpc_mem_121(\PR|prif.pc_mem[12]~13_combout ),
	.imemload_id31(\PR|imemload_id~31_combout ),
	.prifpc_mem_111(\PR|prif.pc_mem[11]~14_combout ),
	.prifpc_mem_101(\PR|prif.pc_mem[10]~15_combout ),
	.prifpc_mem_91(\PR|prif.pc_mem[9]~16_combout ),
	.prifpc_mem_61(\PR|prif.pc_mem[6]~17_combout ),
	.prifpc_mem_271(\PR|prif.pc_mem[27]~18_combout ),
	.prifpc_mem_231(\PR|prif.pc_mem[23]~19_combout ),
	.prifpc_mem_181(\PR|prif.pc_mem[18]~20_combout ),
	.prifpc_mem_241(\PR|prif.pc_mem[24]~21_combout ),
	.prifpc_mem_161(\PR|prif.pc_mem[16]~22_combout ),
	.prifpc_mem_191(\PR|prif.pc_mem[19]~23_combout ),
	.prifpc_mem_171(\PR|prif.pc_mem[17]~24_combout ),
	.prifpc_mem_211(\PR|prif.pc_mem[21]~25_combout ),
	.prifpc_mem_201(\PR|prif.pc_mem[20]~26_combout ),
	.prifpc_mem_261(\PR|prif.pc_mem[26]~27_combout ),
	.prifpc_mem_81(\PR|prif.pc_mem[8]~28_combout ),
	.prifpc_mem_71(\PR|prif.pc_mem[7]~29_combout ),
	.prifpc_mem_221(\PR|prif.pc_mem[22]~30_combout ),
	.prifpc_mem_251(\PR|prif.pc_mem[25]~31_combout ),
	.instr_ex1(\PR|instr_ex~1_combout ),
	.instr_ex2(\PR|instr_ex~2_combout ),
	.instr_ex3(\PR|instr_ex~3_combout ),
	.instr_ex4(\PR|instr_ex~4_combout ),
	.instr_ex5(\PR|instr_ex~5_combout ),
	.instr_ex6(\PR|instr_ex~6_combout ),
	.PCScr_ex(\PR|PCScr_ex~3_combout ),
	.pc_ex(\PR|pc_ex~0_combout ),
	.PCScr_ex1(\PR|PCScr_ex~4_combout ),
	.pc_ex1(\PR|pc_ex~1_combout ),
	.pc_ex2(\PR|pc_ex~2_combout ),
	.pc_ex3(\PR|pc_ex~3_combout ),
	.pc_ex4(\PR|pc_ex~4_combout ),
	.pc_ex5(\PR|pc_ex~5_combout ),
	.pc_ex6(\PR|pc_ex~6_combout ),
	.pc_ex7(\PR|pc_ex~7_combout ),
	.pc_ex8(\PR|pc_ex~8_combout ),
	.pc_ex9(\PR|pc_ex~9_combout ),
	.instr_ex7(\PR|instr_ex~7_combout ),
	.instr_ex8(\PR|instr_ex~8_combout ),
	.pc_ex10(\PR|pc_ex~10_combout ),
	.pc_ex11(\PR|pc_ex~11_combout ),
	.instr_ex9(\PR|instr_ex~9_combout ),
	.instr_ex10(\PR|instr_ex~10_combout ),
	.pc_ex12(\PR|pc_ex~12_combout ),
	.pc_ex13(\PR|pc_ex~13_combout ),
	.instr_ex11(\PR|instr_ex~11_combout ),
	.instr_ex12(\PR|instr_ex~12_combout ),
	.pc_ex14(\PR|pc_ex~14_combout ),
	.pc_ex15(\PR|pc_ex~15_combout ),
	.instr_ex13(\PR|instr_ex~13_combout ),
	.instr_ex14(\PR|instr_ex~14_combout ),
	.pc_ex16(\PR|pc_ex~16_combout ),
	.pc_ex17(\PR|pc_ex~17_combout ),
	.pc_ex18(\PR|pc_ex~18_combout ),
	.pc_ex19(\PR|pc_ex~19_combout ),
	.pc_ex20(\PR|pc_ex~20_combout ),
	.pc_ex21(\PR|pc_ex~21_combout ),
	.pc_ex22(\PR|pc_ex~22_combout ),
	.pc_ex23(\PR|pc_ex~23_combout ),
	.instr_ex15(\PR|instr_ex~15_combout ),
	.instr_ex16(\PR|instr_ex~16_combout ),
	.instr_ex17(\PR|instr_ex~17_combout ),
	.pc_ex24(\PR|pc_ex~24_combout ),
	.pc_ex25(\PR|pc_ex~25_combout ),
	.pc_ex26(\PR|pc_ex~26_combout ),
	.pc_ex27(\PR|pc_ex~27_combout ),
	.pc_ex28(\PR|pc_ex~28_combout ),
	.pc_ex29(\PR|pc_ex~29_combout ),
	.pc_ex30(\PR|pc_ex~30_combout ),
	.pc_ex31(\PR|pc_ex~31_combout ),
	.instr_ex18(\PR|instr_ex~18_combout ),
	.instr_ex19(\PR|instr_ex~19_combout ),
	.instr_ex20(\PR|instr_ex~20_combout ),
	.instr_ex21(\PR|instr_ex~21_combout ),
	.instr_ex22(\PR|instr_ex~22_combout ),
	.instr_ex23(\PR|instr_ex~23_combout ),
	.instr_ex24(\PR|instr_ex~24_combout ),
	.instr_ex25(\PR|instr_ex~25_combout ),
	.halt_wb(\PR|halt_wb~0_combout ),
	.dataScr_ex1(\PR|dataScr_ex~3_combout ),
	.pc_id(\PR|pc_id~0_combout ),
	.pc_id1(\PR|pc_id~1_combout ),
	.pc_id2(\PR|pc_id~2_combout ),
	.pc_id3(\PR|pc_id~3_combout ),
	.pc_id4(\PR|pc_id~4_combout ),
	.pc_id5(\PR|pc_id~5_combout ),
	.pc_id6(\PR|pc_id~6_combout ),
	.pc_id7(\PR|pc_id~7_combout ),
	.pc_id8(\PR|pc_id~8_combout ),
	.pc_id9(\PR|pc_id~9_combout ),
	.pc_id10(\PR|pc_id~10_combout ),
	.pc_id11(\PR|pc_id~11_combout ),
	.pc_id12(\PR|pc_id~12_combout ),
	.pc_id13(\PR|pc_id~13_combout ),
	.pc_id14(\PR|pc_id~14_combout ),
	.pc_id15(\PR|pc_id~15_combout ),
	.pc_id16(\PR|pc_id~16_combout ),
	.pc_id17(\PR|pc_id~17_combout ),
	.pc_id18(\PR|pc_id~18_combout ),
	.pc_id19(\PR|pc_id~19_combout ),
	.pc_id20(\PR|pc_id~20_combout ),
	.pc_id21(\PR|pc_id~21_combout ),
	.pc_id22(\PR|pc_id~22_combout ),
	.pc_id23(\PR|pc_id~23_combout ),
	.pc_id24(\PR|pc_id~24_combout ),
	.pc_id25(\PR|pc_id~25_combout ),
	.pc_id26(\PR|pc_id~26_combout ),
	.pc_id27(\PR|pc_id~27_combout ),
	.pc_id28(\PR|pc_id~28_combout ),
	.pc_id29(\PR|pc_id~29_combout ),
	.pc_id30(\PR|pc_id~30_combout ),
	.pc_id31(\PR|pc_id~31_combout ),
	.dataScr_ex2(\PR|dataScr_ex~4_combout ),
	.ALUScr_ex3(\PR|ALUScr_ex~15_combout ),
	.zero_flag_mem(\PR|zero_flag_mem~13_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

control_unit CU(
	.prifimemload_id_31(\prif.imemload_id [31]),
	.prifimemload_id_30(\prif.imemload_id [30]),
	.prifimemload_id_29(\prif.imemload_id [29]),
	.prifimemload_id_27(\prif.imemload_id [27]),
	.prifimemload_id_26(\prif.imemload_id [26]),
	.prifimemload_id_28(\prif.imemload_id [28]),
	.prifimemload_id_3(\prif.imemload_id [3]),
	.prifimemload_id_1(\prif.imemload_id [1]),
	.prifimemload_id_5(\prif.imemload_id [5]),
	.prifimemload_id_4(\prif.imemload_id [4]),
	.prifimemload_id_2(\prif.imemload_id [2]),
	.prifimemload_id_0(\prif.imemload_id [0]),
	.Equal15(\CU|Equal15~0_combout ),
	.Equal11(\CU|Equal11~0_combout ),
	.Equal0(\CU|Equal0~0_combout ),
	.Equal10(\CU|Equal10~0_combout ),
	.Equal12(\CU|Equal12~0_combout ),
	.Equal20(\CU|Equal20~0_combout ),
	.Equal26(\CU|Equal26~0_combout ),
	.Equal25(\CU|Equal25~1_combout ),
	.Equal13(\CU|Equal13~0_combout ),
	.dataScr_ex(\PR|dataScr_ex~2_combout ),
	.WideNor0(\CU|WideNor0~2_combout ),
	.Selector0(\CU|Selector0~2_combout ),
	.Equal4(\CU|Equal4~0_combout ),
	.Selector2(\CU|Selector2~4_combout ),
	.Selector21(\CU|Selector2~5_combout ),
	.ALUScr_ex(\PR|ALUScr_ex~13_combout ),
	.Selector3(\CU|Selector3~5_combout ),
	.Equal131(\CU|Equal13~1_combout ),
	.ALUScr_ex1(\PR|ALUScr_ex~15_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

alu ALU(
	.prifALUOP_ex_3(\prif.ALUOP_ex [3]),
	.Mux89(\Mux89~2_combout ),
	.Mux94(\Mux94~1_combout ),
	.Mux30(\Mux30~1_combout ),
	.Mux95(\Mux95~1_combout ),
	.Mux31(\Mux31~1_combout ),
	.Mux92(\Mux92~2_combout ),
	.Mux93(\Mux93~0_combout ),
	.Mux61(\Mux61~1_combout ),
	.Mux91(\Mux91~2_combout ),
	.Mux64(\Mux64~0_combout ),
	.Mux65(\Mux65~0_combout ),
	.Mux66(\Mux66~0_combout ),
	.Mux68(\Mux68~0_combout ),
	.Mux72(\Mux72~0_combout ),
	.Mux77(\Mux77~0_combout ),
	.Mux71(\Mux71~0_combout ),
	.Mux79(\Mux79~0_combout ),
	.Mux76(\Mux76~0_combout ),
	.Mux78(\Mux78~0_combout ),
	.Mux74(\Mux74~0_combout ),
	.Mux75(\Mux75~0_combout ),
	.Mux67(\Mux67~0_combout ),
	.Mux69(\Mux69~0_combout ),
	.Mux73(\Mux73~0_combout ),
	.Mux70(\Mux70~0_combout ),
	.prifALUOP_ex_2(\prif.ALUOP_ex [2]),
	.prifALUOP_ex_1(\prif.ALUOP_ex [1]),
	.Mux29(\Mux29~1_combout ),
	.Mux27(\Mux27~1_combout ),
	.Mux28(\Mux28~1_combout ),
	.Mux931(\Mux93~2_combout ),
	.Mux23(\Mux23~1_combout ),
	.Mux24(\Mux24~1_combout ),
	.Mux25(\Mux25~1_combout ),
	.Mux26(\Mux26~1_combout ),
	.Mux15(\Mux15~1_combout ),
	.Mux16(\Mux16~1_combout ),
	.Mux17(\Mux17~1_combout ),
	.Mux18(\Mux18~1_combout ),
	.Mux20(\Mux20~1_combout ),
	.Mux19(\Mux19~0_combout ),
	.Mux191(\Mux19~1_combout ),
	.Mux21(\Mux21~1_combout ),
	.Mux22(\Mux22~1_combout ),
	.Mux13(\Mux13~1_combout ),
	.Mux14(\Mux14~1_combout ),
	.Mux11(\Mux11~1_combout ),
	.Mux12(\Mux12~1_combout ),
	.Mux9(\Mux9~1_combout ),
	.Mux10(\Mux10~1_combout ),
	.Mux7(\Mux7~1_combout ),
	.Mux8(\Mux8~1_combout ),
	.Mux0(\Mux0~1_combout ),
	.Mux1(\Mux1~1_combout ),
	.Mux2(\Mux2~1_combout ),
	.Mux5(\Mux5~1_combout ),
	.Mux6(\Mux6~1_combout ),
	.Mux3(\Mux3~1_combout ),
	.Mux4(\Mux4~1_combout ),
	.prifALUOP_ex_0(\prif.ALUOP_ex [0]),
	.aluifportOut_1(\ALU|aluif.portOut[1]~15_combout ),
	.Mux192(\Mux19~3_combout ),
	.aluifportOut_0(\ALU|aluif.portOut[0]~24_combout ),
	.aluifportOut_3(\ALU|aluif.portOut[3]~30_combout ),
	.aluifportOut_5(\ALU|aluif.portOut[5]~31_combout ),
	.aluifportOut_2(\ALU|aluif.portOut[2]~33_combout ),
	.aluifportOut_31(\ALU|aluif.portOut[3]~39_combout ),
	.aluifportOut_32(\ALU|aluif.portOut[3]~40_combout ),
	.aluifportOut_21(\ALU|aluif.portOut[2]~48_combout ),
	.aluifportOut_51(\ALU|aluif.portOut[5]~57_combout ),
	.aluifportOut_52(\ALU|aluif.portOut[5]~58_combout ),
	.aluifportOut_4(\ALU|aluif.portOut[4]~65_combout ),
	.aluifportOut_7(\ALU|aluif.portOut[7]~72_combout ),
	.aluifportOut_6(\ALU|aluif.portOut[6]~79_combout ),
	.aluifportOut_9(\ALU|aluif.portOut[9]~90_combout ),
	.aluifportOut_8(\ALU|aluif.portOut[8]~96_combout ),
	.aluifportOut_11(\ALU|aluif.portOut[11]~102_combout ),
	.aluifportOut_10(\ALU|aluif.portOut[10]~108_combout ),
	.aluifportOut_13(\ALU|aluif.portOut[13]~114_combout ),
	.aluifportOut_12(\ALU|aluif.portOut[12]~120_combout ),
	.aluifportOut_15(\ALU|aluif.portOut[15]~126_combout ),
	.aluifportOut_14(\ALU|aluif.portOut[14]~132_combout ),
	.aluifportOut_23(\ALU|aluif.portOut[23]~140_combout ),
	.aluifportOut_22(\ALU|aluif.portOut[22]~147_combout ),
	.aluifportOut_211(\ALU|aluif.portOut[21]~153_combout ),
	.aluifportOut_29(\ALU|aluif.portOut[29]~166_combout ),
	.aluifportOut_28(\ALU|aluif.portOut[28]~180_combout ),
	.aluifneg_flag(\ALU|aluif.neg_flag~19_combout ),
	.aluifportOut_30(\ALU|aluif.portOut[30]~189_combout ),
	.aluifportOut_20(\ALU|aluif.portOut[20]~195_combout ),
	.aluifportOut_17(\ALU|aluif.portOut[17]~201_combout ),
	.aluifportOut_16(\ALU|aluif.portOut[16]~207_combout ),
	.aluifportOut_19(\ALU|aluif.portOut[19]~213_combout ),
	.aluifportOut_18(\ALU|aluif.portOut[18]~221_combout ),
	.aluifportOut_25(\ALU|aluif.portOut[25]~234_combout ),
	.aluifportOut_24(\ALU|aluif.portOut[24]~241_combout ),
	.aluifportOut_27(\ALU|aluif.portOut[27]~249_combout ),
	.aluifportOut_26(\ALU|aluif.portOut[26]~257_combout ),
	.aluifportOut_53(\ALU|aluif.portOut[5]~258_combout ),
	.Mux90(\Mux90~3_combout ),
	.Mux80(\Mux80~4_combout ),
	.Mux81(\Mux81~3_combout ),
	.Mux82(\Mux82~3_combout ),
	.Mux83(\Mux83~3_combout ),
	.Mux84(\Mux84~3_combout ),
	.Mux85(\Mux85~3_combout ),
	.Mux86(\Mux86~3_combout ),
	.Mux891(\Mux89~4_combout ),
	.Mux87(\Mux87~3_combout ),
	.Mux88(\Mux88~3_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

register_file RF(
	.prifimemload_id_17(\prif.imemload_id [17]),
	.prifimemload_id_16(\prif.imemload_id [16]),
	.prifimemload_id_19(\prif.imemload_id [19]),
	.prifimemload_id_18(\prif.imemload_id [18]),
	.prifimemload_id_22(\prif.imemload_id [22]),
	.prifimemload_id_21(\prif.imemload_id [21]),
	.prifimemload_id_24(\prif.imemload_id [24]),
	.prifimemload_id_23(\prif.imemload_id [23]),
	.prifRegwen_wb(\prif.Regwen_wb~q ),
	.prifregwrite_wb_2(\prif.regwrite_wb [2]),
	.prifregwrite_wb_0(\prif.regwrite_wb [0]),
	.prifregwrite_wb_1(\prif.regwrite_wb [1]),
	.prifregwrite_wb_4(\prif.regwrite_wb [4]),
	.prifregwrite_wb_3(\prif.regwrite_wb [3]),
	.Equal8(\HU|Equal8~0_combout ),
	.Mux163(\Mux163~1_combout ),
	.Mux164(\Mux164~1_combout ),
	.Mux161(\Mux161~1_combout ),
	.Mux162(\Mux162~1_combout ),
	.Mux160(\Mux160~1_combout ),
	.Mux133(\Mux133~1_combout ),
	.Mux134(\Mux134~1_combout ),
	.Mux135(\Mux135~1_combout ),
	.Mux159(\Mux159~1_combout ),
	.Mux149(\Mux149~1_combout ),
	.Mux150(\Mux150~1_combout ),
	.Mux151(\Mux151~1_combout ),
	.Mux152(\Mux152~1_combout ),
	.Mux153(\Mux153~1_combout ),
	.Mux154(\Mux154~1_combout ),
	.Mux155(\Mux155~1_combout ),
	.Mux158(\Mux158~1_combout ),
	.Mux137(\Mux137~1_combout ),
	.Mux141(\Mux141~1_combout ),
	.Mux146(\Mux146~1_combout ),
	.Mux140(\Mux140~1_combout ),
	.Mux148(\Mux148~1_combout ),
	.Mux145(\Mux145~1_combout ),
	.Mux147(\Mux147~1_combout ),
	.Mux143(\Mux143~1_combout ),
	.Mux144(\Mux144~1_combout ),
	.Mux136(\Mux136~1_combout ),
	.Mux138(\Mux138~1_combout ),
	.Mux156(\Mux156~1_combout ),
	.Mux157(\Mux157~1_combout ),
	.Mux142(\Mux142~1_combout ),
	.Mux139(\Mux139~1_combout ),
	.Mux62(\RF|Mux62~9_combout ),
	.Mux621(\RF|Mux62~19_combout ),
	.Mux30(\RF|Mux30~9_combout ),
	.Mux301(\RF|Mux30~19_combout ),
	.Mux63(\RF|Mux63~9_combout ),
	.Mux631(\RF|Mux63~19_combout ),
	.Mux31(\RF|Mux31~9_combout ),
	.Mux311(\RF|Mux31~19_combout ),
	.Mux60(\RF|Mux60~9_combout ),
	.Mux601(\RF|Mux60~19_combout ),
	.Mux61(\RF|Mux61~9_combout ),
	.Mux611(\RF|Mux61~19_combout ),
	.Mux59(\RF|Mux59~9_combout ),
	.Mux591(\RF|Mux59~19_combout ),
	.Mux32(\RF|Mux32~9_combout ),
	.Mux321(\RF|Mux32~19_combout ),
	.Mux33(\RF|Mux33~9_combout ),
	.Mux331(\RF|Mux33~19_combout ),
	.Mux34(\RF|Mux34~9_combout ),
	.Mux341(\RF|Mux34~19_combout ),
	.Mux58(\RF|Mux58~9_combout ),
	.Mux581(\RF|Mux58~19_combout ),
	.Mux48(\RF|Mux48~9_combout ),
	.Mux481(\RF|Mux48~19_combout ),
	.Mux49(\RF|Mux49~9_combout ),
	.Mux491(\RF|Mux49~19_combout ),
	.Mux50(\RF|Mux50~9_combout ),
	.Mux501(\RF|Mux50~19_combout ),
	.Mux51(\RF|Mux51~9_combout ),
	.Mux511(\RF|Mux51~19_combout ),
	.Mux52(\RF|Mux52~9_combout ),
	.Mux521(\RF|Mux52~19_combout ),
	.Mux53(\RF|Mux53~9_combout ),
	.Mux531(\RF|Mux53~19_combout ),
	.Mux54(\RF|Mux54~9_combout ),
	.Mux541(\RF|Mux54~19_combout ),
	.Mux57(\RF|Mux57~9_combout ),
	.Mux571(\RF|Mux57~19_combout ),
	.Mux36(\RF|Mux36~9_combout ),
	.Mux361(\RF|Mux36~19_combout ),
	.Mux40(\RF|Mux40~9_combout ),
	.Mux401(\RF|Mux40~19_combout ),
	.Mux45(\RF|Mux45~9_combout ),
	.Mux451(\RF|Mux45~19_combout ),
	.Mux39(\RF|Mux39~9_combout ),
	.Mux391(\RF|Mux39~19_combout ),
	.Mux47(\RF|Mux47~9_combout ),
	.Mux471(\RF|Mux47~19_combout ),
	.Mux44(\RF|Mux44~9_combout ),
	.Mux441(\RF|Mux44~19_combout ),
	.Mux46(\RF|Mux46~9_combout ),
	.Mux461(\RF|Mux46~19_combout ),
	.Mux42(\RF|Mux42~9_combout ),
	.Mux421(\RF|Mux42~19_combout ),
	.Mux43(\RF|Mux43~9_combout ),
	.Mux431(\RF|Mux43~19_combout ),
	.Mux35(\RF|Mux35~9_combout ),
	.Mux351(\RF|Mux35~19_combout ),
	.Mux37(\RF|Mux37~9_combout ),
	.Mux371(\RF|Mux37~19_combout ),
	.Mux55(\RF|Mux55~9_combout ),
	.Mux551(\RF|Mux55~19_combout ),
	.Mux56(\RF|Mux56~9_combout ),
	.Mux561(\RF|Mux56~19_combout ),
	.Mux41(\RF|Mux41~9_combout ),
	.Mux411(\RF|Mux41~19_combout ),
	.Mux38(\RF|Mux38~9_combout ),
	.Mux381(\RF|Mux38~19_combout ),
	.Mux29(\RF|Mux29~9_combout ),
	.Mux291(\RF|Mux29~19_combout ),
	.Mux27(\RF|Mux27~9_combout ),
	.Mux271(\RF|Mux27~19_combout ),
	.Mux28(\RF|Mux28~9_combout ),
	.Mux281(\RF|Mux28~19_combout ),
	.Mux23(\RF|Mux23~9_combout ),
	.Mux231(\RF|Mux23~19_combout ),
	.Mux24(\RF|Mux24~9_combout ),
	.Mux241(\RF|Mux24~19_combout ),
	.Mux25(\RF|Mux25~9_combout ),
	.Mux251(\RF|Mux25~19_combout ),
	.Mux26(\RF|Mux26~9_combout ),
	.Mux261(\RF|Mux26~19_combout ),
	.Mux15(\RF|Mux15~9_combout ),
	.Mux1510(\RF|Mux15~19_combout ),
	.Mux16(\RF|Mux16~9_combout ),
	.Mux165(\RF|Mux16~19_combout ),
	.Mux17(\RF|Mux17~9_combout ),
	.Mux171(\RF|Mux17~19_combout ),
	.Mux18(\RF|Mux18~9_combout ),
	.Mux181(\RF|Mux18~19_combout ),
	.Mux20(\RF|Mux20~9_combout ),
	.Mux201(\RF|Mux20~19_combout ),
	.Mux19(\RF|Mux19~9_combout ),
	.Mux191(\RF|Mux19~19_combout ),
	.Mux21(\RF|Mux21~9_combout ),
	.Mux211(\RF|Mux21~19_combout ),
	.Mux22(\RF|Mux22~9_combout ),
	.Mux221(\RF|Mux22~19_combout ),
	.Mux13(\RF|Mux13~9_combout ),
	.Mux131(\RF|Mux13~19_combout ),
	.Mux14(\RF|Mux14~9_combout ),
	.Mux1410(\RF|Mux14~19_combout ),
	.Mux11(\RF|Mux11~9_combout ),
	.Mux111(\RF|Mux11~19_combout ),
	.Mux12(\RF|Mux12~9_combout ),
	.Mux121(\RF|Mux12~19_combout ),
	.Mux9(\RF|Mux9~9_combout ),
	.Mux91(\RF|Mux9~19_combout ),
	.Mux10(\RF|Mux10~9_combout ),
	.Mux101(\RF|Mux10~19_combout ),
	.Mux7(\RF|Mux7~9_combout ),
	.Mux71(\RF|Mux7~19_combout ),
	.Mux8(\RF|Mux8~9_combout ),
	.Mux81(\RF|Mux8~19_combout ),
	.Mux0(\RF|Mux0~9_combout ),
	.Mux01(\RF|Mux0~19_combout ),
	.Mux1(\RF|Mux1~9_combout ),
	.Mux110(\RF|Mux1~19_combout ),
	.Mux2(\RF|Mux2~9_combout ),
	.Mux210(\RF|Mux2~19_combout ),
	.Mux5(\RF|Mux5~9_combout ),
	.Mux510(\RF|Mux5~19_combout ),
	.Mux6(\RF|Mux6~9_combout ),
	.Mux64(\RF|Mux6~19_combout ),
	.Mux3(\RF|Mux3~9_combout ),
	.Mux310(\RF|Mux3~19_combout ),
	.Mux4(\RF|Mux4~9_combout ),
	.Mux410(\RF|Mux4~19_combout ),
	.CLK(CLK),
	.nRST(nRST1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X55_Y23_N29
dffeas \prif.imm_ex[1] (
	.clk(CLK),
	.d(\PR|imm_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[1] .is_wysiwyg = "true";
defparam \prif.imm_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N5
dffeas \prif.ALUScr_ex[1] (
	.clk(CLK),
	.d(\PR|ALUScr_ex~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.ALUScr_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.ALUScr_ex[1] .is_wysiwyg = "true";
defparam \prif.ALUScr_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y23_N31
dffeas \prif.shamt_ex[1] (
	.clk(CLK),
	.d(\PR|shamt_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.shamt_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.shamt_ex[1] .is_wysiwyg = "true";
defparam \prif.shamt_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N5
dffeas \prif.ALUScr_ex[0] (
	.clk(CLK),
	.d(\prif.ALUScr_ex[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.ALUScr_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.ALUScr_ex[0] .is_wysiwyg = "true";
defparam \prif.ALUScr_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N13
dffeas \prif.Regwen_mem (
	.clk(CLK),
	.d(\PR|Regwen_mem~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.Regwen_mem~q ),
	.prn(vcc));
// synopsys translate_off
defparam \prif.Regwen_mem .is_wysiwyg = "true";
defparam \prif.Regwen_mem .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N11
dffeas \prif.regwrite_mem[4] (
	.clk(CLK),
	.d(\PR|regwrite_mem~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_mem [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_mem[4] .is_wysiwyg = "true";
defparam \prif.regwrite_mem[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N5
dffeas \prif.regwrite_mem[0] (
	.clk(CLK),
	.d(\PR|regwrite_mem~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_mem [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_mem[0] .is_wysiwyg = "true";
defparam \prif.regwrite_mem[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N27
dffeas \prif.regwrite_mem[1] (
	.clk(CLK),
	.d(\PR|regwrite_mem~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_mem [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_mem[1] .is_wysiwyg = "true";
defparam \prif.regwrite_mem[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N1
dffeas \prif.regwrite_mem[2] (
	.clk(CLK),
	.d(\PR|regwrite_mem~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_mem [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_mem[2] .is_wysiwyg = "true";
defparam \prif.regwrite_mem[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N23
dffeas \prif.regwrite_mem[3] (
	.clk(CLK),
	.d(\PR|regwrite_mem~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_mem [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_mem[3] .is_wysiwyg = "true";
defparam \prif.regwrite_mem[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y27_N25
dffeas \prif.rt_ex[1] (
	.clk(CLK),
	.d(\PR|rt_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rt_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rt_ex[1] .is_wysiwyg = "true";
defparam \prif.rt_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y27_N3
dffeas \prif.rt_ex[0] (
	.clk(CLK),
	.d(\PR|rt_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rt_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rt_ex[0] .is_wysiwyg = "true";
defparam \prif.rt_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y27_N5
dffeas \prif.rt_ex[3] (
	.clk(CLK),
	.d(\PR|rt_ex~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rt_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rt_ex[3] .is_wysiwyg = "true";
defparam \prif.rt_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y27_N11
dffeas \prif.rt_ex[2] (
	.clk(CLK),
	.d(\PR|rt_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rt_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rt_ex[2] .is_wysiwyg = "true";
defparam \prif.rt_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y27_N9
dffeas \prif.rt_ex[4] (
	.clk(CLK),
	.d(\PR|rt_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rt_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rt_ex[4] .is_wysiwyg = "true";
defparam \prif.rt_ex[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y27_N21
dffeas \prif.rdat2_ex[1] (
	.clk(CLK),
	.d(\PR|rdat2_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[1] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N1
dffeas \prif.opcode_mem[1] (
	.clk(CLK),
	.d(\PR|opcode_mem~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_mem [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_mem[1] .is_wysiwyg = "true";
defparam \prif.opcode_mem[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N7
dffeas \prif.opcode_mem[0] (
	.clk(CLK),
	.d(\PR|opcode_mem~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_mem [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_mem[0] .is_wysiwyg = "true";
defparam \prif.opcode_mem[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N13
dffeas \prif.opcode_mem[2] (
	.clk(CLK),
	.d(\PR|opcode_mem~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_mem [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_mem[2] .is_wysiwyg = "true";
defparam \prif.opcode_mem[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N3
dffeas \prif.opcode_mem[3] (
	.clk(CLK),
	.d(\PR|opcode_mem~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_mem [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_mem[3] .is_wysiwyg = "true";
defparam \prif.opcode_mem[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N25
dffeas \prif.opcode_mem[5] (
	.clk(CLK),
	.d(\PR|opcode_mem~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_mem [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_mem[5] .is_wysiwyg = "true";
defparam \prif.opcode_mem[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y30_N27
dffeas \prif.opcode_mem[4] (
	.clk(CLK),
	.d(\PR|opcode_mem~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_mem [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_mem[4] .is_wysiwyg = "true";
defparam \prif.opcode_mem[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y25_N29
dffeas \prif.rdat1_ex[1] (
	.clk(CLK),
	.d(\PR|rdat1_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[1] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N9
dffeas \prif.imm_ex[0] (
	.clk(CLK),
	.d(\PR|imm_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[0] .is_wysiwyg = "true";
defparam \prif.imm_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N3
dffeas \prif.shamt_ex[0] (
	.clk(CLK),
	.d(\PR|shamt_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.shamt_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.shamt_ex[0] .is_wysiwyg = "true";
defparam \prif.shamt_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N17
dffeas \prif.rdat2_ex[0] (
	.clk(CLK),
	.d(\PR|rdat2_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[0] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y25_N11
dffeas \prif.rdat1_ex[0] (
	.clk(CLK),
	.d(\PR|rdat1_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[0] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N1
dffeas \prif.rdat2_ex[3] (
	.clk(CLK),
	.d(\PR|rdat2_ex~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[3] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N19
dffeas \prif.imm_ex[3] (
	.clk(CLK),
	.d(\PR|imm_ex~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[3] .is_wysiwyg = "true";
defparam \prif.imm_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y28_N29
dffeas \prif.shamt_ex[3] (
	.clk(CLK),
	.d(\PR|shamt_ex~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.shamt_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.shamt_ex[3] .is_wysiwyg = "true";
defparam \prif.shamt_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N13
dffeas \prif.imm_ex[2] (
	.clk(CLK),
	.d(\PR|imm_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[2] .is_wysiwyg = "true";
defparam \prif.imm_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y23_N21
dffeas \prif.shamt_ex[2] (
	.clk(CLK),
	.d(\PR|shamt_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.shamt_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.shamt_ex[2] .is_wysiwyg = "true";
defparam \prif.shamt_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N23
dffeas \prif.rdat2_ex[2] (
	.clk(CLK),
	.d(\PR|rdat2_ex~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[2] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y27_N31
dffeas \prif.rdat2_ex[4] (
	.clk(CLK),
	.d(\PR|rdat2_ex~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[4] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N27
dffeas \prif.imm_ex[4] (
	.clk(CLK),
	.d(\PR|imm_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[4] .is_wysiwyg = "true";
defparam \prif.imm_ex[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N5
dffeas \prif.shamt_ex[4] (
	.clk(CLK),
	.d(\PR|shamt_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.shamt_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.shamt_ex[4] .is_wysiwyg = "true";
defparam \prif.shamt_ex[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N21
dffeas \prif.instr_ex[15] (
	.clk(CLK),
	.d(\PR|instr_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[15] .is_wysiwyg = "true";
defparam \prif.instr_ex[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y25_N5
dffeas \prif.rdat2_ex[31] (
	.clk(CLK),
	.d(\PR|rdat2_ex~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[31] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N23
dffeas \prif.imm_mem[15] (
	.clk(CLK),
	.d(\PR|imm_mem~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[15] .is_wysiwyg = "true";
defparam \prif.imm_mem[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y27_N1
dffeas \prif.rdat2_ex[30] (
	.clk(CLK),
	.d(\PR|rdat2_ex~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[30] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N27
dffeas \prif.imm_mem[14] (
	.clk(CLK),
	.d(\PR|imm_mem~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[14] .is_wysiwyg = "true";
defparam \prif.imm_mem[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y27_N7
dffeas \prif.rdat2_ex[29] (
	.clk(CLK),
	.d(\PR|rdat2_ex~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[29] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N3
dffeas \prif.imm_mem[13] (
	.clk(CLK),
	.d(\PR|imm_mem~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[13] .is_wysiwyg = "true";
defparam \prif.imm_mem[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N17
dffeas \prif.imm_ex[5] (
	.clk(CLK),
	.d(\PR|imm_ex~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[5] .is_wysiwyg = "true";
defparam \prif.imm_ex[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N5
dffeas \prif.rdat2_ex[5] (
	.clk(CLK),
	.d(\PR|rdat2_ex~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[5] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N23
dffeas \prif.imm_ex[15] (
	.clk(CLK),
	.d(\PR|imm_ex~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[15] .is_wysiwyg = "true";
defparam \prif.imm_ex[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y27_N29
dffeas \prif.rdat2_ex[15] (
	.clk(CLK),
	.d(\PR|rdat2_ex~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[15] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N17
dffeas \prif.imm_ex[14] (
	.clk(CLK),
	.d(\PR|imm_ex~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[14] .is_wysiwyg = "true";
defparam \prif.imm_ex[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N21
dffeas \prif.rdat2_ex[14] (
	.clk(CLK),
	.d(\PR|rdat2_ex~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[14] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y26_N29
dffeas \prif.imm_ex[13] (
	.clk(CLK),
	.d(\PR|imm_ex~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[13] .is_wysiwyg = "true";
defparam \prif.imm_ex[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y26_N27
dffeas \prif.rdat2_ex[13] (
	.clk(CLK),
	.d(\PR|rdat2_ex~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[13] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N1
dffeas \prif.imm_ex[12] (
	.clk(CLK),
	.d(\PR|imm_ex~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[12] .is_wysiwyg = "true";
defparam \prif.imm_ex[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N11
dffeas \prif.rdat2_ex[12] (
	.clk(CLK),
	.d(\PR|rdat2_ex~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[12] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y27_N23
dffeas \prif.imm_ex[11] (
	.clk(CLK),
	.d(\PR|imm_ex~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[11] .is_wysiwyg = "true";
defparam \prif.imm_ex[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N27
dffeas \prif.rdat2_ex[11] (
	.clk(CLK),
	.d(\PR|rdat2_ex~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[11] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N11
dffeas \prif.imm_ex[10] (
	.clk(CLK),
	.d(\PR|imm_ex~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[10] .is_wysiwyg = "true";
defparam \prif.imm_ex[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y26_N1
dffeas \prif.rdat2_ex[10] (
	.clk(CLK),
	.d(\PR|rdat2_ex~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[10] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N11
dffeas \prif.imm_ex[9] (
	.clk(CLK),
	.d(\PR|imm_ex~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[9] .is_wysiwyg = "true";
defparam \prif.imm_ex[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N5
dffeas \prif.rdat2_ex[9] (
	.clk(CLK),
	.d(\PR|rdat2_ex~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[9] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N5
dffeas \prif.imm_ex[6] (
	.clk(CLK),
	.d(\PR|imm_ex~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[6] .is_wysiwyg = "true";
defparam \prif.imm_ex[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N31
dffeas \prif.rdat2_ex[6] (
	.clk(CLK),
	.d(\PR|rdat2_ex~33_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[6] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N21
dffeas \prif.rdat2_ex[27] (
	.clk(CLK),
	.d(\PR|rdat2_ex~35_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[27] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y26_N31
dffeas \prif.imm_mem[11] (
	.clk(CLK),
	.d(\PR|imm_mem~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[11] .is_wysiwyg = "true";
defparam \prif.imm_mem[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N27
dffeas \prif.rdat2_ex[23] (
	.clk(CLK),
	.d(\PR|rdat2_ex~37_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[23] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N17
dffeas \prif.imm_mem[7] (
	.clk(CLK),
	.d(\PR|imm_mem~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[7] .is_wysiwyg = "true";
defparam \prif.imm_mem[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N9
dffeas \prif.rdat2_ex[18] (
	.clk(CLK),
	.d(\PR|rdat2_ex~39_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[18] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N9
dffeas \prif.imm_mem[2] (
	.clk(CLK),
	.d(\PR|imm_mem~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[2] .is_wysiwyg = "true";
defparam \prif.imm_mem[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N19
dffeas \prif.rdat2_ex[24] (
	.clk(CLK),
	.d(\PR|rdat2_ex~41_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[24] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N13
dffeas \prif.imm_mem[8] (
	.clk(CLK),
	.d(\PR|imm_mem~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[8] .is_wysiwyg = "true";
defparam \prif.imm_mem[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N5
dffeas \prif.rdat2_ex[16] (
	.clk(CLK),
	.d(\PR|rdat2_ex~43_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[16] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N3
dffeas \prif.imm_mem[0] (
	.clk(CLK),
	.d(\PR|imm_mem~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[0] .is_wysiwyg = "true";
defparam \prif.imm_mem[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N27
dffeas \prif.rdat2_ex[19] (
	.clk(CLK),
	.d(\PR|rdat2_ex~45_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[19] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N27
dffeas \prif.imm_mem[3] (
	.clk(CLK),
	.d(\PR|imm_mem~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[3] .is_wysiwyg = "true";
defparam \prif.imm_mem[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y27_N9
dffeas \prif.rdat2_ex[17] (
	.clk(CLK),
	.d(\PR|rdat2_ex~47_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[17] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N29
dffeas \prif.imm_mem[1] (
	.clk(CLK),
	.d(\PR|imm_mem~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[1] .is_wysiwyg = "true";
defparam \prif.imm_mem[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N21
dffeas \prif.rdat2_ex[21] (
	.clk(CLK),
	.d(\PR|rdat2_ex~49_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[21] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N5
dffeas \prif.imm_mem[5] (
	.clk(CLK),
	.d(\PR|imm_mem~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[5] .is_wysiwyg = "true";
defparam \prif.imm_mem[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N5
dffeas \prif.rdat2_ex[20] (
	.clk(CLK),
	.d(\PR|rdat2_ex~51_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[20] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N31
dffeas \prif.imm_mem[4] (
	.clk(CLK),
	.d(\PR|imm_mem~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[4] .is_wysiwyg = "true";
defparam \prif.imm_mem[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N25
dffeas \prif.rdat2_ex[28] (
	.clk(CLK),
	.d(\PR|rdat2_ex~53_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[28] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y26_N9
dffeas \prif.imm_mem[12] (
	.clk(CLK),
	.d(\PR|imm_mem~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[12] .is_wysiwyg = "true";
defparam \prif.imm_mem[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N9
dffeas \prif.rdat2_ex[26] (
	.clk(CLK),
	.d(\PR|rdat2_ex~55_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[26] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N27
dffeas \prif.imm_mem[10] (
	.clk(CLK),
	.d(\PR|imm_mem~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[10] .is_wysiwyg = "true";
defparam \prif.imm_mem[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N15
dffeas \prif.imm_ex[8] (
	.clk(CLK),
	.d(\PR|imm_ex~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[8] .is_wysiwyg = "true";
defparam \prif.imm_ex[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N31
dffeas \prif.rdat2_ex[8] (
	.clk(CLK),
	.d(\PR|rdat2_ex~57_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[8] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y23_N11
dffeas \prif.imm_ex[7] (
	.clk(CLK),
	.d(\PR|imm_ex~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_ex [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_ex[7] .is_wysiwyg = "true";
defparam \prif.imm_ex[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N17
dffeas \prif.rdat2_ex[7] (
	.clk(CLK),
	.d(\PR|rdat2_ex~59_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[7] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y27_N13
dffeas \prif.rdat2_ex[22] (
	.clk(CLK),
	.d(\PR|rdat2_ex~61_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[22] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y26_N1
dffeas \prif.imm_mem[6] (
	.clk(CLK),
	.d(\PR|imm_mem~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[6] .is_wysiwyg = "true";
defparam \prif.imm_mem[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N25
dffeas \prif.rdat2_ex[25] (
	.clk(CLK),
	.d(\PR|rdat2_ex~63_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat2_ex [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat2_ex[25] .is_wysiwyg = "true";
defparam \prif.rdat2_ex[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N25
dffeas \prif.imm_mem[9] (
	.clk(CLK),
	.d(\PR|imm_mem~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_mem [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_mem[9] .is_wysiwyg = "true";
defparam \prif.imm_mem[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y25_N9
dffeas \prif.rdat1_ex[2] (
	.clk(CLK),
	.d(\PR|rdat1_ex~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[2] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N1
dffeas \prif.rdat1_ex[4] (
	.clk(CLK),
	.d(\PR|rdat1_ex~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[4] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N31
dffeas \prif.rdat1_ex[3] (
	.clk(CLK),
	.d(\PR|rdat1_ex~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[3] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N31
dffeas \prif.rdat1_ex[8] (
	.clk(CLK),
	.d(\PR|rdat1_ex~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[8] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y25_N31
dffeas \prif.rdat1_ex[7] (
	.clk(CLK),
	.d(\PR|rdat1_ex~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[7] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N1
dffeas \prif.rdat1_ex[6] (
	.clk(CLK),
	.d(\PR|rdat1_ex~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[6] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N5
dffeas \prif.rdat1_ex[5] (
	.clk(CLK),
	.d(\PR|rdat1_ex~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[5] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N23
dffeas \prif.rdat1_ex[16] (
	.clk(CLK),
	.d(\PR|rdat1_ex~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[16] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N15
dffeas \prif.rdat1_ex[15] (
	.clk(CLK),
	.d(\PR|rdat1_ex~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[15] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N29
dffeas \prif.rdat1_ex[14] (
	.clk(CLK),
	.d(\PR|rdat1_ex~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[14] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y26_N21
dffeas \prif.rdat1_ex[13] (
	.clk(CLK),
	.d(\PR|rdat1_ex~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[13] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N23
dffeas \prif.rdat1_ex[11] (
	.clk(CLK),
	.d(\PR|rdat1_ex~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[11] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N13
dffeas \prif.rdat1_ex[12] (
	.clk(CLK),
	.d(\PR|rdat1_ex~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[12] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N23
dffeas \prif.rdat1_ex[10] (
	.clk(CLK),
	.d(\PR|rdat1_ex~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[10] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y26_N27
dffeas \prif.rdat1_ex[9] (
	.clk(CLK),
	.d(\PR|rdat1_ex~33_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[9] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N29
dffeas \prif.rdat1_ex[18] (
	.clk(CLK),
	.d(\PR|rdat1_ex~35_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[18] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N15
dffeas \prif.rdat1_ex[17] (
	.clk(CLK),
	.d(\PR|rdat1_ex~37_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[17] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N7
dffeas \prif.rdat1_ex[20] (
	.clk(CLK),
	.d(\PR|rdat1_ex~39_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[20] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y26_N9
dffeas \prif.rdat1_ex[19] (
	.clk(CLK),
	.d(\PR|rdat1_ex~41_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[19] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N29
dffeas \prif.rdat1_ex[22] (
	.clk(CLK),
	.d(\PR|rdat1_ex~43_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[22] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N15
dffeas \prif.rdat1_ex[21] (
	.clk(CLK),
	.d(\PR|rdat1_ex~45_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[21] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N13
dffeas \prif.rdat1_ex[24] (
	.clk(CLK),
	.d(\PR|rdat1_ex~47_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[24] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N3
dffeas \prif.rdat1_ex[23] (
	.clk(CLK),
	.d(\PR|rdat1_ex~49_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[23] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N1
dffeas \prif.rdat1_ex[31] (
	.clk(CLK),
	.d(\PR|rdat1_ex~51_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[31] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N27
dffeas \prif.rdat1_ex[30] (
	.clk(CLK),
	.d(\PR|rdat1_ex~53_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[30] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y34_N25
dffeas \prif.rdat1_ex[29] (
	.clk(CLK),
	.d(\PR|rdat1_ex~55_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[29] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N25
dffeas \prif.rdat1_ex[26] (
	.clk(CLK),
	.d(\PR|rdat1_ex~57_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[26] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N15
dffeas \prif.rdat1_ex[25] (
	.clk(CLK),
	.d(\PR|rdat1_ex~59_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[25] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N5
dffeas \prif.rdat1_ex[28] (
	.clk(CLK),
	.d(\PR|rdat1_ex~61_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[28] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y34_N23
dffeas \prif.rdat1_ex[27] (
	.clk(CLK),
	.d(\PR|rdat1_ex~63_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_ex [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_ex[27] .is_wysiwyg = "true";
defparam \prif.rdat1_ex[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N29
dffeas \prif.opcode_ex[5] (
	.clk(CLK),
	.d(\PR|opcode_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_ex [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_ex[5] .is_wysiwyg = "true";
defparam \prif.opcode_ex[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N5
dffeas \prif.opcode_ex[0] (
	.clk(CLK),
	.d(\PR|opcode_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_ex[0] .is_wysiwyg = "true";
defparam \prif.opcode_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N15
dffeas \prif.opcode_ex[1] (
	.clk(CLK),
	.d(\PR|opcode_ex~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_ex[1] .is_wysiwyg = "true";
defparam \prif.opcode_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N5
dffeas \prif.opcode_ex[2] (
	.clk(CLK),
	.d(\PR|opcode_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_ex[2] .is_wysiwyg = "true";
defparam \prif.opcode_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N29
dffeas \prif.opcode_ex[4] (
	.clk(CLK),
	.d(\PR|opcode_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_ex[4] .is_wysiwyg = "true";
defparam \prif.opcode_ex[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N13
dffeas \prif.memren_ex (
	.clk(CLK),
	.d(\PR|memren_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.memren_ex~q ),
	.prn(vcc));
// synopsys translate_off
defparam \prif.memren_ex .is_wysiwyg = "true";
defparam \prif.memren_ex .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N27
dffeas \prif.memwen_ex (
	.clk(CLK),
	.d(\PR|memwen_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.memwen_ex~q ),
	.prn(vcc));
// synopsys translate_off
defparam \prif.memwen_ex .is_wysiwyg = "true";
defparam \prif.memwen_ex .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N5
dffeas \prif.pc_bran_mem[3] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[3] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y33_N1
dffeas \prif.pc_bran_mem[4] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[4] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N16
cycloneive_lcell_comb \Add3~14 (
// Equation(s):
// \Add3~14_combout  = (pc_9 & (!\Add3~13 )) # (!pc_9 & ((\Add3~13 ) # (GND)))
// \Add3~15  = CARRY((!\Add3~13 ) # (!pc_9))

	.dataa(pc_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~13 ),
	.combout(\Add3~14_combout ),
	.cout(\Add3~15 ));
// synopsys translate_off
defparam \Add3~14 .lut_mask = 16'h5A5F;
defparam \Add3~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X56_Y33_N27
dffeas \prif.rdat1_mem[8] (
	.clk(CLK),
	.d(\PR|rdat1_mem~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[8] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y28_N19
dffeas \prif.rdat1_mem[10] (
	.clk(CLK),
	.d(\PR|rdat1_mem~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[10] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N0
cycloneive_lcell_comb \Add3~30 (
// Equation(s):
// \Add3~30_combout  = (pc_17 & (!\Add3~29 )) # (!pc_17 & ((\Add3~29 ) # (GND)))
// \Add3~31  = CARRY((!\Add3~29 ) # (!pc_17))

	.dataa(pc_17),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~29 ),
	.combout(\Add3~30_combout ),
	.cout(\Add3~31 ));
// synopsys translate_off
defparam \Add3~30 .lut_mask = 16'h5A5F;
defparam \Add3~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N4
cycloneive_lcell_comb \Add3~34 (
// Equation(s):
// \Add3~34_combout  = (pc_19 & (!\Add3~33 )) # (!pc_19 & ((\Add3~33 ) # (GND)))
// \Add3~35  = CARRY((!\Add3~33 ) # (!pc_19))

	.dataa(pc_19),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~33 ),
	.combout(\Add3~34_combout ),
	.cout(\Add3~35 ));
// synopsys translate_off
defparam \Add3~34 .lut_mask = 16'h5A5F;
defparam \Add3~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X57_Y30_N31
dffeas \prif.pc_bran_mem[23] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[23] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N11
dffeas \prif.pc_bran_mem[22] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[22] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N16
cycloneive_lcell_comb \Add3~46 (
// Equation(s):
// \Add3~46_combout  = (pc_25 & (!\Add3~45 )) # (!pc_25 & ((\Add3~45 ) # (GND)))
// \Add3~47  = CARRY((!\Add3~45 ) # (!pc_25))

	.dataa(pc_25),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~45 ),
	.combout(\Add3~46_combout ),
	.cout(\Add3~47 ));
// synopsys translate_off
defparam \Add3~46 .lut_mask = 16'h5A5F;
defparam \Add3~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X55_Y32_N31
dffeas \prif.pc_bran_mem[29] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[29] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N23
dffeas \prif.pc_bran_mem[20] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[20] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N15
dffeas \prif.halt_ex (
	.clk(CLK),
	.d(\PR|halt_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.halt_ex~q ),
	.prn(vcc));
// synopsys translate_off
defparam \prif.halt_ex .is_wysiwyg = "true";
defparam \prif.halt_ex .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N21
dffeas \prif.imemload_id[31] (
	.clk(CLK),
	.d(\PR|imemload_id~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[31] .is_wysiwyg = "true";
defparam \prif.imemload_id[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N23
dffeas \prif.imemload_id[30] (
	.clk(CLK),
	.d(\PR|imemload_id~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[30] .is_wysiwyg = "true";
defparam \prif.imemload_id[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N25
dffeas \prif.imemload_id[29] (
	.clk(CLK),
	.d(\PR|imemload_id~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[29] .is_wysiwyg = "true";
defparam \prif.imemload_id[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N15
dffeas \prif.imemload_id[27] (
	.clk(CLK),
	.d(\PR|imemload_id~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[27] .is_wysiwyg = "true";
defparam \prif.imemload_id[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N17
dffeas \prif.imemload_id[26] (
	.clk(CLK),
	.d(\PR|imemload_id~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[26] .is_wysiwyg = "true";
defparam \prif.imemload_id[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N7
dffeas \prif.imemload_id[28] (
	.clk(CLK),
	.d(\PR|imemload_id~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[28] .is_wysiwyg = "true";
defparam \prif.imemload_id[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y27_N25
dffeas \prif.imemload_id[3] (
	.clk(CLK),
	.d(\PR|imemload_id~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[3] .is_wysiwyg = "true";
defparam \prif.imemload_id[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y28_N9
dffeas \prif.imemload_id[1] (
	.clk(CLK),
	.d(\PR|imemload_id~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[1] .is_wysiwyg = "true";
defparam \prif.imemload_id[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y27_N27
dffeas \prif.imemload_id[5] (
	.clk(CLK),
	.d(\PR|imemload_id~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[5] .is_wysiwyg = "true";
defparam \prif.imemload_id[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y27_N29
dffeas \prif.imemload_id[4] (
	.clk(CLK),
	.d(\PR|imemload_id~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[4] .is_wysiwyg = "true";
defparam \prif.imemload_id[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y27_N15
dffeas \prif.imemload_id[2] (
	.clk(CLK),
	.d(\PR|imemload_id~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[2] .is_wysiwyg = "true";
defparam \prif.imemload_id[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y27_N17
dffeas \prif.imemload_id[0] (
	.clk(CLK),
	.d(\PR|imemload_id~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[0] .is_wysiwyg = "true";
defparam \prif.imemload_id[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y28_N31
dffeas \prif.imemload_id[7] (
	.clk(CLK),
	.d(\PR|imemload_id~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[7] .is_wysiwyg = "true";
defparam \prif.imemload_id[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N7
dffeas \prif.Regwen_ex (
	.clk(CLK),
	.d(\PR|Regwen_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.Regwen_ex~q ),
	.prn(vcc));
// synopsys translate_off
defparam \prif.Regwen_ex .is_wysiwyg = "true";
defparam \prif.Regwen_ex .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N25
dffeas \prif.rd_ex[4] (
	.clk(CLK),
	.d(\PR|rd_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rd_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rd_ex[4] .is_wysiwyg = "true";
defparam \prif.rd_ex[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N13
dffeas \prif.RegDest_ex[1] (
	.clk(CLK),
	.d(\PR|RegDest_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.RegDest_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.RegDest_ex[1] .is_wysiwyg = "true";
defparam \prif.RegDest_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N19
dffeas \prif.RegDest_ex[0] (
	.clk(CLK),
	.d(\PR|RegDest_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.RegDest_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.RegDest_ex[0] .is_wysiwyg = "true";
defparam \prif.RegDest_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y27_N19
dffeas \prif.rd_ex[0] (
	.clk(CLK),
	.d(\PR|rd_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rd_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rd_ex[0] .is_wysiwyg = "true";
defparam \prif.rd_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N29
dffeas \prif.rd_ex[1] (
	.clk(CLK),
	.d(\PR|rd_ex~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rd_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rd_ex[1] .is_wysiwyg = "true";
defparam \prif.rd_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N7
dffeas \prif.rd_ex[2] (
	.clk(CLK),
	.d(\PR|rd_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rd_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rd_ex[2] .is_wysiwyg = "true";
defparam \prif.rd_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N3
dffeas \prif.rd_ex[3] (
	.clk(CLK),
	.d(\PR|rd_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rd_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rd_ex[3] .is_wysiwyg = "true";
defparam \prif.rd_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N9
dffeas \prif.imemload_id[17] (
	.clk(CLK),
	.d(\PR|imemload_id~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[17] .is_wysiwyg = "true";
defparam \prif.imemload_id[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N15
dffeas \prif.imemload_id[16] (
	.clk(CLK),
	.d(\PR|imemload_id~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[16] .is_wysiwyg = "true";
defparam \prif.imemload_id[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N9
dffeas \prif.imemload_id[19] (
	.clk(CLK),
	.d(\PR|imemload_id~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[19] .is_wysiwyg = "true";
defparam \prif.imemload_id[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N1
dffeas \prif.imemload_id[18] (
	.clk(CLK),
	.d(\PR|imemload_id~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[18] .is_wysiwyg = "true";
defparam \prif.imemload_id[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y31_N5
dffeas \prif.imemload_id[20] (
	.clk(CLK),
	.d(\PR|imemload_id~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[20] .is_wysiwyg = "true";
defparam \prif.imemload_id[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N1
dffeas \prif.dataScr_mem[0] (
	.clk(CLK),
	.d(\PR|dataScr_mem~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dataScr_mem [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dataScr_mem[0] .is_wysiwyg = "true";
defparam \prif.dataScr_mem[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N29
dffeas \prif.dataScr_mem[1] (
	.clk(CLK),
	.d(\PR|dataScr_mem~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dataScr_mem [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dataScr_mem[1] .is_wysiwyg = "true";
defparam \prif.dataScr_mem[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N29
dffeas \prif.imemload_id[22] (
	.clk(CLK),
	.d(\PR|imemload_id~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[22] .is_wysiwyg = "true";
defparam \prif.imemload_id[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N27
dffeas \prif.imemload_id[21] (
	.clk(CLK),
	.d(\PR|imemload_id~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[21] .is_wysiwyg = "true";
defparam \prif.imemload_id[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N3
dffeas \prif.imemload_id[24] (
	.clk(CLK),
	.d(\PR|imemload_id~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[24] .is_wysiwyg = "true";
defparam \prif.imemload_id[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N1
dffeas \prif.imemload_id[23] (
	.clk(CLK),
	.d(\PR|imemload_id~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[23] .is_wysiwyg = "true";
defparam \prif.imemload_id[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y28_N13
dffeas \prif.imemload_id[25] (
	.clk(CLK),
	.d(\PR|imemload_id~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[25] .is_wysiwyg = "true";
defparam \prif.imemload_id[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N13
dffeas \prif.opcode_ex[3] (
	.clk(CLK),
	.d(\PR|opcode_ex~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.opcode_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.opcode_ex[3] .is_wysiwyg = "true";
defparam \prif.opcode_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y28_N19
dffeas \prif.imemload_id[6] (
	.clk(CLK),
	.d(\PR|imemload_id~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[6] .is_wysiwyg = "true";
defparam \prif.imemload_id[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y28_N5
dffeas \prif.imemload_id[9] (
	.clk(CLK),
	.d(\PR|imemload_id~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[9] .is_wysiwyg = "true";
defparam \prif.imemload_id[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N25
dffeas \prif.imemload_id[8] (
	.clk(CLK),
	.d(\PR|imemload_id~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[8] .is_wysiwyg = "true";
defparam \prif.imemload_id[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N3
dffeas \prif.imemload_id[10] (
	.clk(CLK),
	.d(\PR|imemload_id~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[10] .is_wysiwyg = "true";
defparam \prif.imemload_id[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N19
dffeas \prif.imemload_id[15] (
	.clk(CLK),
	.d(\PR|imemload_id~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[15] .is_wysiwyg = "true";
defparam \prif.imemload_id[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N5
dffeas \prif.imemload_id[14] (
	.clk(CLK),
	.d(\PR|imemload_id~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[14] .is_wysiwyg = "true";
defparam \prif.imemload_id[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N5
dffeas \prif.imemload_id[13] (
	.clk(CLK),
	.d(\PR|imemload_id~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[13] .is_wysiwyg = "true";
defparam \prif.imemload_id[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y32_N27
dffeas \prif.imemload_id[12] (
	.clk(CLK),
	.d(\PR|imemload_id~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[12] .is_wysiwyg = "true";
defparam \prif.imemload_id[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N19
dffeas \prif.imemload_id[11] (
	.clk(CLK),
	.d(\PR|imemload_id~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imemload_id [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imemload_id[11] .is_wysiwyg = "true";
defparam \prif.imemload_id[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N31
dffeas \prif.instr_ex[3] (
	.clk(CLK),
	.d(\PR|instr_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[3] .is_wysiwyg = "true";
defparam \prif.instr_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N11
dffeas \prif.instr_ex[5] (
	.clk(CLK),
	.d(\PR|instr_ex~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[5] .is_wysiwyg = "true";
defparam \prif.instr_ex[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N29
dffeas \prif.instr_ex[4] (
	.clk(CLK),
	.d(\PR|instr_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[4] .is_wysiwyg = "true";
defparam \prif.instr_ex[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N7
dffeas \prif.instr_ex[2] (
	.clk(CLK),
	.d(\PR|instr_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[2] .is_wysiwyg = "true";
defparam \prif.instr_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y23_N1
dffeas \prif.instr_ex[1] (
	.clk(CLK),
	.d(\PR|instr_ex~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[1] .is_wysiwyg = "true";
defparam \prif.instr_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N3
dffeas \prif.instr_ex[0] (
	.clk(CLK),
	.d(\PR|instr_ex~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[0] .is_wysiwyg = "true";
defparam \prif.instr_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y32_N29
dffeas \prif.PCScr_ex[0] (
	.clk(CLK),
	.d(\PR|PCScr_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.PCScr_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.PCScr_ex[0] .is_wysiwyg = "true";
defparam \prif.PCScr_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N31
dffeas \prif.pc_ex[1] (
	.clk(CLK),
	.d(\PR|pc_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[1] .is_wysiwyg = "true";
defparam \prif.pc_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N5
dffeas \prif.PCScr_ex[1] (
	.clk(CLK),
	.d(\PR|PCScr_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.PCScr_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.PCScr_ex[1] .is_wysiwyg = "true";
defparam \prif.PCScr_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N17
dffeas \prif.pc_ex[0] (
	.clk(CLK),
	.d(\PR|pc_ex~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[0] .is_wysiwyg = "true";
defparam \prif.pc_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N21
dffeas \prif.pc_ex[3] (
	.clk(CLK),
	.d(\PR|pc_ex~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[3] .is_wysiwyg = "true";
defparam \prif.pc_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N9
dffeas \prif.pc_ex[2] (
	.clk(CLK),
	.d(\PR|pc_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[2] .is_wysiwyg = "true";
defparam \prif.pc_ex[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N2
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (\prif.pc_ex [2] & (\prif.imm_ex [0] $ (VCC))) # (!\prif.pc_ex [2] & (\prif.imm_ex [0] & VCC))
// \Add0~1  = CARRY((\prif.pc_ex [2] & \prif.imm_ex [0]))

	.dataa(\prif.pc_ex [2]),
	.datab(\prif.imm_ex [0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h6688;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N4
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (\prif.imm_ex [1] & ((\prif.pc_ex [3] & (\Add0~1  & VCC)) # (!\prif.pc_ex [3] & (!\Add0~1 )))) # (!\prif.imm_ex [1] & ((\prif.pc_ex [3] & (!\Add0~1 )) # (!\prif.pc_ex [3] & ((\Add0~1 ) # (GND)))))
// \Add0~3  = CARRY((\prif.imm_ex [1] & (!\prif.pc_ex [3] & !\Add0~1 )) # (!\prif.imm_ex [1] & ((!\Add0~1 ) # (!\prif.pc_ex [3]))))

	.dataa(\prif.imm_ex [1]),
	.datab(\prif.pc_ex [3]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h9617;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X56_Y32_N1
dffeas \prif.pc_ex[5] (
	.clk(CLK),
	.d(\PR|pc_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[5] .is_wysiwyg = "true";
defparam \prif.pc_ex[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N23
dffeas \prif.pc_ex[4] (
	.clk(CLK),
	.d(\PR|pc_ex~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[4] .is_wysiwyg = "true";
defparam \prif.pc_ex[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N6
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = ((\prif.pc_ex [4] $ (\prif.imm_ex [2] $ (!\Add0~3 )))) # (GND)
// \Add0~5  = CARRY((\prif.pc_ex [4] & ((\prif.imm_ex [2]) # (!\Add0~3 ))) # (!\prif.pc_ex [4] & (\prif.imm_ex [2] & !\Add0~3 )))

	.dataa(\prif.pc_ex [4]),
	.datab(\prif.imm_ex [2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h698E;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N8
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (\prif.imm_ex [3] & ((\prif.pc_ex [5] & (\Add0~5  & VCC)) # (!\prif.pc_ex [5] & (!\Add0~5 )))) # (!\prif.imm_ex [3] & ((\prif.pc_ex [5] & (!\Add0~5 )) # (!\prif.pc_ex [5] & ((\Add0~5 ) # (GND)))))
// \Add0~7  = CARRY((\prif.imm_ex [3] & (!\prif.pc_ex [5] & !\Add0~5 )) # (!\prif.imm_ex [3] & ((!\Add0~5 ) # (!\prif.pc_ex [5]))))

	.dataa(\prif.imm_ex [3]),
	.datab(\prif.pc_ex [5]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h9617;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X54_Y33_N31
dffeas \prif.pc_ex[7] (
	.clk(CLK),
	.d(\PR|pc_ex~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[7] .is_wysiwyg = "true";
defparam \prif.pc_ex[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N13
dffeas \prif.pc_ex[6] (
	.clk(CLK),
	.d(\PR|pc_ex~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[6] .is_wysiwyg = "true";
defparam \prif.pc_ex[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N10
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = ((\prif.pc_ex [6] $ (\prif.imm_ex [4] $ (!\Add0~7 )))) # (GND)
// \Add0~9  = CARRY((\prif.pc_ex [6] & ((\prif.imm_ex [4]) # (!\Add0~7 ))) # (!\prif.pc_ex [6] & (\prif.imm_ex [4] & !\Add0~7 )))

	.dataa(\prif.pc_ex [6]),
	.datab(\prif.imm_ex [4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h698E;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N12
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (\prif.imm_ex [5] & ((\prif.pc_ex [7] & (\Add0~9  & VCC)) # (!\prif.pc_ex [7] & (!\Add0~9 )))) # (!\prif.imm_ex [5] & ((\prif.pc_ex [7] & (!\Add0~9 )) # (!\prif.pc_ex [7] & ((\Add0~9 ) # (GND)))))
// \Add0~11  = CARRY((\prif.imm_ex [5] & (!\prif.pc_ex [7] & !\Add0~9 )) # (!\prif.imm_ex [5] & ((!\Add0~9 ) # (!\prif.pc_ex [7]))))

	.dataa(\prif.imm_ex [5]),
	.datab(\prif.pc_ex [7]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h9617;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X54_Y33_N11
dffeas \prif.pc_ex[9] (
	.clk(CLK),
	.d(\PR|pc_ex~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[9] .is_wysiwyg = "true";
defparam \prif.pc_ex[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N17
dffeas \prif.pc_ex[8] (
	.clk(CLK),
	.d(\PR|pc_ex~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[8] .is_wysiwyg = "true";
defparam \prif.pc_ex[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N14
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = ((\prif.pc_ex [8] $ (\prif.imm_ex [6] $ (!\Add0~11 )))) # (GND)
// \Add0~13  = CARRY((\prif.pc_ex [8] & ((\prif.imm_ex [6]) # (!\Add0~11 ))) # (!\prif.pc_ex [8] & (\prif.imm_ex [6] & !\Add0~11 )))

	.dataa(\prif.pc_ex [8]),
	.datab(\prif.imm_ex [6]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h698E;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N16
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (\prif.pc_ex [9] & ((\prif.imm_ex [7] & (\Add0~13  & VCC)) # (!\prif.imm_ex [7] & (!\Add0~13 )))) # (!\prif.pc_ex [9] & ((\prif.imm_ex [7] & (!\Add0~13 )) # (!\prif.imm_ex [7] & ((\Add0~13 ) # (GND)))))
// \Add0~15  = CARRY((\prif.pc_ex [9] & (!\prif.imm_ex [7] & !\Add0~13 )) # (!\prif.pc_ex [9] & ((!\Add0~13 ) # (!\prif.imm_ex [7]))))

	.dataa(\prif.pc_ex [9]),
	.datab(\prif.imm_ex [7]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h9617;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X55_Y23_N7
dffeas \prif.instr_ex[7] (
	.clk(CLK),
	.d(\PR|instr_ex~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[7] .is_wysiwyg = "true";
defparam \prif.instr_ex[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N7
dffeas \prif.instr_ex[6] (
	.clk(CLK),
	.d(\PR|instr_ex~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[6] .is_wysiwyg = "true";
defparam \prif.instr_ex[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N29
dffeas \prif.pc_ex[11] (
	.clk(CLK),
	.d(\PR|pc_ex~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[11] .is_wysiwyg = "true";
defparam \prif.pc_ex[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N3
dffeas \prif.pc_ex[10] (
	.clk(CLK),
	.d(\PR|pc_ex~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[10] .is_wysiwyg = "true";
defparam \prif.pc_ex[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N18
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = ((\prif.imm_ex [8] $ (\prif.pc_ex [10] $ (!\Add0~15 )))) # (GND)
// \Add0~17  = CARRY((\prif.imm_ex [8] & ((\prif.pc_ex [10]) # (!\Add0~15 ))) # (!\prif.imm_ex [8] & (\prif.pc_ex [10] & !\Add0~15 )))

	.dataa(\prif.imm_ex [8]),
	.datab(\prif.pc_ex [10]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N20
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (\prif.imm_ex [9] & ((\prif.pc_ex [11] & (\Add0~17  & VCC)) # (!\prif.pc_ex [11] & (!\Add0~17 )))) # (!\prif.imm_ex [9] & ((\prif.pc_ex [11] & (!\Add0~17 )) # (!\prif.pc_ex [11] & ((\Add0~17 ) # (GND)))))
// \Add0~19  = CARRY((\prif.imm_ex [9] & (!\prif.pc_ex [11] & !\Add0~17 )) # (!\prif.imm_ex [9] & ((!\Add0~17 ) # (!\prif.pc_ex [11]))))

	.dataa(\prif.imm_ex [9]),
	.datab(\prif.pc_ex [11]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h9617;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X61_Y32_N9
dffeas \prif.instr_ex[9] (
	.clk(CLK),
	.d(\PR|instr_ex~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[9] .is_wysiwyg = "true";
defparam \prif.instr_ex[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N13
dffeas \prif.instr_ex[8] (
	.clk(CLK),
	.d(\PR|instr_ex~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[8] .is_wysiwyg = "true";
defparam \prif.instr_ex[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N1
dffeas \prif.pc_ex[13] (
	.clk(CLK),
	.d(\PR|pc_ex~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[13] .is_wysiwyg = "true";
defparam \prif.pc_ex[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N19
dffeas \prif.pc_ex[12] (
	.clk(CLK),
	.d(\PR|pc_ex~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[12] .is_wysiwyg = "true";
defparam \prif.pc_ex[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N22
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = ((\prif.imm_ex [10] $ (\prif.pc_ex [12] $ (!\Add0~19 )))) # (GND)
// \Add0~21  = CARRY((\prif.imm_ex [10] & ((\prif.pc_ex [12]) # (!\Add0~19 ))) # (!\prif.imm_ex [10] & (\prif.pc_ex [12] & !\Add0~19 )))

	.dataa(\prif.imm_ex [10]),
	.datab(\prif.pc_ex [12]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h698E;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N24
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (\prif.pc_ex [13] & ((\prif.imm_ex [11] & (\Add0~21  & VCC)) # (!\prif.imm_ex [11] & (!\Add0~21 )))) # (!\prif.pc_ex [13] & ((\prif.imm_ex [11] & (!\Add0~21 )) # (!\prif.imm_ex [11] & ((\Add0~21 ) # (GND)))))
// \Add0~23  = CARRY((\prif.pc_ex [13] & (!\prif.imm_ex [11] & !\Add0~21 )) # (!\prif.pc_ex [13] & ((!\Add0~21 ) # (!\prif.imm_ex [11]))))

	.dataa(\prif.pc_ex [13]),
	.datab(\prif.imm_ex [11]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h9617;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X54_Y27_N25
dffeas \prif.instr_ex[11] (
	.clk(CLK),
	.d(\PR|instr_ex~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[11] .is_wysiwyg = "true";
defparam \prif.instr_ex[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N15
dffeas \prif.instr_ex[10] (
	.clk(CLK),
	.d(\PR|instr_ex~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[10] .is_wysiwyg = "true";
defparam \prif.instr_ex[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N21
dffeas \prif.pc_ex[15] (
	.clk(CLK),
	.d(\PR|pc_ex~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[15] .is_wysiwyg = "true";
defparam \prif.pc_ex[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N31
dffeas \prif.pc_ex[14] (
	.clk(CLK),
	.d(\PR|pc_ex~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[14] .is_wysiwyg = "true";
defparam \prif.pc_ex[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N26
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = ((\prif.pc_ex [14] $ (\prif.imm_ex [12] $ (!\Add0~23 )))) # (GND)
// \Add0~25  = CARRY((\prif.pc_ex [14] & ((\prif.imm_ex [12]) # (!\Add0~23 ))) # (!\prif.pc_ex [14] & (\prif.imm_ex [12] & !\Add0~23 )))

	.dataa(\prif.pc_ex [14]),
	.datab(\prif.imm_ex [12]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'h698E;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N28
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (\prif.pc_ex [15] & ((\prif.imm_ex [13] & (\Add0~25  & VCC)) # (!\prif.imm_ex [13] & (!\Add0~25 )))) # (!\prif.pc_ex [15] & ((\prif.imm_ex [13] & (!\Add0~25 )) # (!\prif.imm_ex [13] & ((\Add0~25 ) # (GND)))))
// \Add0~27  = CARRY((\prif.pc_ex [15] & (!\prif.imm_ex [13] & !\Add0~25 )) # (!\prif.pc_ex [15] & ((!\Add0~25 ) # (!\prif.imm_ex [13]))))

	.dataa(\prif.pc_ex [15]),
	.datab(\prif.imm_ex [13]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h9617;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X57_Y33_N11
dffeas \prif.instr_ex[13] (
	.clk(CLK),
	.d(\PR|instr_ex~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[13] .is_wysiwyg = "true";
defparam \prif.instr_ex[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N15
dffeas \prif.instr_ex[12] (
	.clk(CLK),
	.d(\PR|instr_ex~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[12] .is_wysiwyg = "true";
defparam \prif.instr_ex[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N11
dffeas \prif.pc_ex[23] (
	.clk(CLK),
	.d(\PR|pc_ex~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[23] .is_wysiwyg = "true";
defparam \prif.pc_ex[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N9
dffeas \prif.pc_ex[22] (
	.clk(CLK),
	.d(\PR|pc_ex~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[22] .is_wysiwyg = "true";
defparam \prif.pc_ex[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N1
dffeas \prif.pc_ex[21] (
	.clk(CLK),
	.d(\PR|pc_ex~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[21] .is_wysiwyg = "true";
defparam \prif.pc_ex[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N1
dffeas \prif.pc_ex[20] (
	.clk(CLK),
	.d(\PR|pc_ex~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[20] .is_wysiwyg = "true";
defparam \prif.pc_ex[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N3
dffeas \prif.pc_ex[19] (
	.clk(CLK),
	.d(\PR|pc_ex~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[19] .is_wysiwyg = "true";
defparam \prif.pc_ex[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N13
dffeas \prif.pc_ex[18] (
	.clk(CLK),
	.d(\PR|pc_ex~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[18] .is_wysiwyg = "true";
defparam \prif.pc_ex[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N27
dffeas \prif.pc_ex[17] (
	.clk(CLK),
	.d(\PR|pc_ex~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[17] .is_wysiwyg = "true";
defparam \prif.pc_ex[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N9
dffeas \prif.pc_ex[16] (
	.clk(CLK),
	.d(\PR|pc_ex~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[16] .is_wysiwyg = "true";
defparam \prif.pc_ex[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N30
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = ((\prif.imm_ex [14] $ (\prif.pc_ex [16] $ (!\Add0~27 )))) # (GND)
// \Add0~29  = CARRY((\prif.imm_ex [14] & ((\prif.pc_ex [16]) # (!\Add0~27 ))) # (!\prif.imm_ex [14] & (\prif.pc_ex [16] & !\Add0~27 )))

	.dataa(\prif.imm_ex [14]),
	.datab(\prif.pc_ex [16]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'h698E;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N0
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (\prif.pc_ex [17] & ((\prif.imm_ex [15] & (\Add0~29  & VCC)) # (!\prif.imm_ex [15] & (!\Add0~29 )))) # (!\prif.pc_ex [17] & ((\prif.imm_ex [15] & (!\Add0~29 )) # (!\prif.imm_ex [15] & ((\Add0~29 ) # (GND)))))
// \Add0~31  = CARRY((\prif.pc_ex [17] & (!\prif.imm_ex [15] & !\Add0~29 )) # (!\prif.pc_ex [17] & ((!\Add0~29 ) # (!\prif.imm_ex [15]))))

	.dataa(\prif.pc_ex [17]),
	.datab(\prif.imm_ex [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h9617;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N2
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = ((\prif.pc_ex [18] $ (\prif.imm_ex [15] $ (!\Add0~31 )))) # (GND)
// \Add0~33  = CARRY((\prif.pc_ex [18] & ((\prif.imm_ex [15]) # (!\Add0~31 ))) # (!\prif.pc_ex [18] & (\prif.imm_ex [15] & !\Add0~31 )))

	.dataa(\prif.pc_ex [18]),
	.datab(\prif.imm_ex [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'h698E;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N4
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (\prif.pc_ex [19] & ((\prif.imm_ex [15] & (\Add0~33  & VCC)) # (!\prif.imm_ex [15] & (!\Add0~33 )))) # (!\prif.pc_ex [19] & ((\prif.imm_ex [15] & (!\Add0~33 )) # (!\prif.imm_ex [15] & ((\Add0~33 ) # (GND)))))
// \Add0~35  = CARRY((\prif.pc_ex [19] & (!\prif.imm_ex [15] & !\Add0~33 )) # (!\prif.pc_ex [19] & ((!\Add0~33 ) # (!\prif.imm_ex [15]))))

	.dataa(\prif.pc_ex [19]),
	.datab(\prif.imm_ex [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h9617;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N6
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = ((\prif.pc_ex [20] $ (\prif.imm_ex [15] $ (!\Add0~35 )))) # (GND)
// \Add0~37  = CARRY((\prif.pc_ex [20] & ((\prif.imm_ex [15]) # (!\Add0~35 ))) # (!\prif.pc_ex [20] & (\prif.imm_ex [15] & !\Add0~35 )))

	.dataa(\prif.pc_ex [20]),
	.datab(\prif.imm_ex [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'h698E;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N8
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (\prif.pc_ex [21] & ((\prif.imm_ex [15] & (\Add0~37  & VCC)) # (!\prif.imm_ex [15] & (!\Add0~37 )))) # (!\prif.pc_ex [21] & ((\prif.imm_ex [15] & (!\Add0~37 )) # (!\prif.imm_ex [15] & ((\Add0~37 ) # (GND)))))
// \Add0~39  = CARRY((\prif.pc_ex [21] & (!\prif.imm_ex [15] & !\Add0~37 )) # (!\prif.pc_ex [21] & ((!\Add0~37 ) # (!\prif.imm_ex [15]))))

	.dataa(\prif.pc_ex [21]),
	.datab(\prif.imm_ex [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h9617;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N10
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = ((\prif.pc_ex [22] $ (\prif.imm_ex [15] $ (!\Add0~39 )))) # (GND)
// \Add0~41  = CARRY((\prif.pc_ex [22] & ((\prif.imm_ex [15]) # (!\Add0~39 ))) # (!\prif.pc_ex [22] & (\prif.imm_ex [15] & !\Add0~39 )))

	.dataa(\prif.pc_ex [22]),
	.datab(\prif.imm_ex [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'h698E;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N12
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// \Add0~42_combout  = (\prif.imm_ex [15] & ((\prif.pc_ex [23] & (\Add0~41  & VCC)) # (!\prif.pc_ex [23] & (!\Add0~41 )))) # (!\prif.imm_ex [15] & ((\prif.pc_ex [23] & (!\Add0~41 )) # (!\prif.pc_ex [23] & ((\Add0~41 ) # (GND)))))
// \Add0~43  = CARRY((\prif.imm_ex [15] & (!\prif.pc_ex [23] & !\Add0~41 )) # (!\prif.imm_ex [15] & ((!\Add0~41 ) # (!\prif.pc_ex [23]))))

	.dataa(\prif.imm_ex [15]),
	.datab(\prif.pc_ex [23]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(\Add0~42_combout ),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h9617;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X55_Y31_N31
dffeas \prif.instr_ex[21] (
	.clk(CLK),
	.d(\PR|instr_ex~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[21] .is_wysiwyg = "true";
defparam \prif.instr_ex[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N21
dffeas \prif.instr_ex[20] (
	.clk(CLK),
	.d(\PR|instr_ex~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[20] .is_wysiwyg = "true";
defparam \prif.instr_ex[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N17
dffeas \prif.instr_ex[19] (
	.clk(CLK),
	.d(\PR|instr_ex~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[19] .is_wysiwyg = "true";
defparam \prif.instr_ex[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N15
dffeas \prif.pc_ex[29] (
	.clk(CLK),
	.d(\PR|pc_ex~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[29] .is_wysiwyg = "true";
defparam \prif.pc_ex[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N3
dffeas \prif.pc_ex[28] (
	.clk(CLK),
	.d(\PR|pc_ex~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[28] .is_wysiwyg = "true";
defparam \prif.pc_ex[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N11
dffeas \prif.pc_ex[27] (
	.clk(CLK),
	.d(\PR|pc_ex~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[27] .is_wysiwyg = "true";
defparam \prif.pc_ex[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N25
dffeas \prif.pc_ex[26] (
	.clk(CLK),
	.d(\PR|pc_ex~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[26] .is_wysiwyg = "true";
defparam \prif.pc_ex[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N13
dffeas \prif.pc_ex[25] (
	.clk(CLK),
	.d(\PR|pc_ex~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[25] .is_wysiwyg = "true";
defparam \prif.pc_ex[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N5
dffeas \prif.pc_ex[24] (
	.clk(CLK),
	.d(\PR|pc_ex~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[24] .is_wysiwyg = "true";
defparam \prif.pc_ex[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N14
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// \Add0~44_combout  = ((\prif.pc_ex [24] $ (\prif.imm_ex [15] $ (!\Add0~43 )))) # (GND)
// \Add0~45  = CARRY((\prif.pc_ex [24] & ((\prif.imm_ex [15]) # (!\Add0~43 ))) # (!\prif.pc_ex [24] & (\prif.imm_ex [15] & !\Add0~43 )))

	.dataa(\prif.pc_ex [24]),
	.datab(\prif.imm_ex [15]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(\Add0~44_combout ),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'h698E;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N16
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = (\prif.imm_ex [15] & ((\prif.pc_ex [25] & (\Add0~45  & VCC)) # (!\prif.pc_ex [25] & (!\Add0~45 )))) # (!\prif.imm_ex [15] & ((\prif.pc_ex [25] & (!\Add0~45 )) # (!\prif.pc_ex [25] & ((\Add0~45 ) # (GND)))))
// \Add0~47  = CARRY((\prif.imm_ex [15] & (!\prif.pc_ex [25] & !\Add0~45 )) # (!\prif.imm_ex [15] & ((!\Add0~45 ) # (!\prif.pc_ex [25]))))

	.dataa(\prif.imm_ex [15]),
	.datab(\prif.pc_ex [25]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(\Add0~46_combout ),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h9617;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N18
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// \Add0~48_combout  = ((\prif.imm_ex [15] $ (\prif.pc_ex [26] $ (!\Add0~47 )))) # (GND)
// \Add0~49  = CARRY((\prif.imm_ex [15] & ((\prif.pc_ex [26]) # (!\Add0~47 ))) # (!\prif.imm_ex [15] & (\prif.pc_ex [26] & !\Add0~47 )))

	.dataa(\prif.imm_ex [15]),
	.datab(\prif.pc_ex [26]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(\Add0~48_combout ),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'h698E;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N20
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// \Add0~50_combout  = (\prif.imm_ex [15] & ((\prif.pc_ex [27] & (\Add0~49  & VCC)) # (!\prif.pc_ex [27] & (!\Add0~49 )))) # (!\prif.imm_ex [15] & ((\prif.pc_ex [27] & (!\Add0~49 )) # (!\prif.pc_ex [27] & ((\Add0~49 ) # (GND)))))
// \Add0~51  = CARRY((\prif.imm_ex [15] & (!\prif.pc_ex [27] & !\Add0~49 )) # (!\prif.imm_ex [15] & ((!\Add0~49 ) # (!\prif.pc_ex [27]))))

	.dataa(\prif.imm_ex [15]),
	.datab(\prif.pc_ex [27]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(\Add0~50_combout ),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h9617;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N22
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = ((\prif.imm_ex [15] $ (\prif.pc_ex [28] $ (!\Add0~51 )))) # (GND)
// \Add0~53  = CARRY((\prif.imm_ex [15] & ((\prif.pc_ex [28]) # (!\Add0~51 ))) # (!\prif.imm_ex [15] & (\prif.pc_ex [28] & !\Add0~51 )))

	.dataa(\prif.imm_ex [15]),
	.datab(\prif.pc_ex [28]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(\Add0~52_combout ),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'h698E;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N24
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// \Add0~54_combout  = (\prif.imm_ex [15] & ((\prif.pc_ex [29] & (\Add0~53  & VCC)) # (!\prif.pc_ex [29] & (!\Add0~53 )))) # (!\prif.imm_ex [15] & ((\prif.pc_ex [29] & (!\Add0~53 )) # (!\prif.pc_ex [29] & ((\Add0~53 ) # (GND)))))
// \Add0~55  = CARRY((\prif.imm_ex [15] & (!\prif.pc_ex [29] & !\Add0~53 )) # (!\prif.imm_ex [15] & ((!\Add0~53 ) # (!\prif.pc_ex [29]))))

	.dataa(\prif.imm_ex [15]),
	.datab(\prif.pc_ex [29]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(\Add0~54_combout ),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h9617;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X55_Y34_N1
dffeas \prif.pc_ex[31] (
	.clk(CLK),
	.d(\PR|pc_ex~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[31] .is_wysiwyg = "true";
defparam \prif.pc_ex[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N15
dffeas \prif.pc_ex[30] (
	.clk(CLK),
	.d(\PR|pc_ex~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_ex [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_ex[30] .is_wysiwyg = "true";
defparam \prif.pc_ex[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N26
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// \Add0~56_combout  = ((\prif.imm_ex [15] $ (\prif.pc_ex [30] $ (!\Add0~55 )))) # (GND)
// \Add0~57  = CARRY((\prif.imm_ex [15] & ((\prif.pc_ex [30]) # (!\Add0~55 ))) # (!\prif.imm_ex [15] & (\prif.pc_ex [30] & !\Add0~55 )))

	.dataa(\prif.imm_ex [15]),
	.datab(\prif.pc_ex [30]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(\Add0~56_combout ),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'h698E;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N28
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = \prif.pc_ex [31] $ (\Add0~57  $ (\prif.imm_ex [15]))

	.dataa(gnd),
	.datab(\prif.pc_ex [31]),
	.datac(gnd),
	.datad(\prif.imm_ex [15]),
	.cin(\Add0~57 ),
	.combout(\Add0~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'hC33C;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X61_Y32_N31
dffeas \prif.instr_ex[18] (
	.clk(CLK),
	.d(\PR|instr_ex~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[18] .is_wysiwyg = "true";
defparam \prif.instr_ex[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N31
dffeas \prif.instr_ex[14] (
	.clk(CLK),
	.d(\PR|instr_ex~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[14] .is_wysiwyg = "true";
defparam \prif.instr_ex[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N31
dffeas \prif.instr_ex[17] (
	.clk(CLK),
	.d(\PR|instr_ex~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[17] .is_wysiwyg = "true";
defparam \prif.instr_ex[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N17
dffeas \prif.instr_ex[16] (
	.clk(CLK),
	.d(\PR|instr_ex~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[16] .is_wysiwyg = "true";
defparam \prif.instr_ex[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y32_N3
dffeas \prif.instr_ex[23] (
	.clk(CLK),
	.d(\PR|instr_ex~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[23] .is_wysiwyg = "true";
defparam \prif.instr_ex[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N25
dffeas \prif.instr_ex[22] (
	.clk(CLK),
	.d(\PR|instr_ex~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[22] .is_wysiwyg = "true";
defparam \prif.instr_ex[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N9
dffeas \prif.instr_ex[25] (
	.clk(CLK),
	.d(\PR|instr_ex~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[25] .is_wysiwyg = "true";
defparam \prif.instr_ex[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N29
dffeas \prif.instr_ex[24] (
	.clk(CLK),
	.d(\PR|instr_ex~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_ex [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_ex[24] .is_wysiwyg = "true";
defparam \prif.instr_ex[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N31
dffeas \prif.dataScr_ex[0] (
	.clk(CLK),
	.d(\PR|dataScr_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dataScr_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dataScr_ex[0] .is_wysiwyg = "true";
defparam \prif.dataScr_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N21
dffeas \prif.dataScr_ex[1] (
	.clk(CLK),
	.d(\PR|dataScr_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|flush_idex~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dataScr_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dataScr_ex[1] .is_wysiwyg = "true";
defparam \prif.dataScr_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N9
dffeas \prif.pc_id[1] (
	.clk(CLK),
	.d(\PR|pc_id~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[1] .is_wysiwyg = "true";
defparam \prif.pc_id[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N7
dffeas \prif.pc_id[0] (
	.clk(CLK),
	.d(\PR|pc_id~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[0] .is_wysiwyg = "true";
defparam \prif.pc_id[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N5
dffeas \prif.pc_id[3] (
	.clk(CLK),
	.d(\PR|pc_id~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[3] .is_wysiwyg = "true";
defparam \prif.pc_id[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N17
dffeas \prif.pc_id[2] (
	.clk(CLK),
	.d(\PR|pc_id~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[2] .is_wysiwyg = "true";
defparam \prif.pc_id[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N23
dffeas \prif.pc_id[5] (
	.clk(CLK),
	.d(\PR|pc_id~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[5] .is_wysiwyg = "true";
defparam \prif.pc_id[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N7
dffeas \prif.pc_id[4] (
	.clk(CLK),
	.d(\PR|pc_id~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[4] .is_wysiwyg = "true";
defparam \prif.pc_id[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N5
dffeas \prif.pc_id[7] (
	.clk(CLK),
	.d(\PR|pc_id~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[7] .is_wysiwyg = "true";
defparam \prif.pc_id[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N31
dffeas \prif.pc_id[6] (
	.clk(CLK),
	.d(\PR|pc_id~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[6] .is_wysiwyg = "true";
defparam \prif.pc_id[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N21
dffeas \prif.pc_id[9] (
	.clk(CLK),
	.d(\PR|pc_id~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[9] .is_wysiwyg = "true";
defparam \prif.pc_id[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N19
dffeas \prif.pc_id[8] (
	.clk(CLK),
	.d(\PR|pc_id~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[8] .is_wysiwyg = "true";
defparam \prif.pc_id[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N1
dffeas \prif.pc_id[11] (
	.clk(CLK),
	.d(\PR|pc_id~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[11] .is_wysiwyg = "true";
defparam \prif.pc_id[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N13
dffeas \prif.pc_id[10] (
	.clk(CLK),
	.d(\PR|pc_id~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[10] .is_wysiwyg = "true";
defparam \prif.pc_id[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N29
dffeas \prif.pc_id[13] (
	.clk(CLK),
	.d(\PR|pc_id~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[13] .is_wysiwyg = "true";
defparam \prif.pc_id[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y33_N3
dffeas \prif.pc_id[12] (
	.clk(CLK),
	.d(\PR|pc_id~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[12] .is_wysiwyg = "true";
defparam \prif.pc_id[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N31
dffeas \prif.pc_id[15] (
	.clk(CLK),
	.d(\PR|pc_id~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[15] .is_wysiwyg = "true";
defparam \prif.pc_id[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N11
dffeas \prif.pc_id[14] (
	.clk(CLK),
	.d(\PR|pc_id~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[14] .is_wysiwyg = "true";
defparam \prif.pc_id[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y32_N31
dffeas \prif.pc_id[23] (
	.clk(CLK),
	.d(\PR|pc_id~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[23] .is_wysiwyg = "true";
defparam \prif.pc_id[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N13
dffeas \prif.pc_id[22] (
	.clk(CLK),
	.d(\PR|pc_id~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[22] .is_wysiwyg = "true";
defparam \prif.pc_id[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N25
dffeas \prif.pc_id[21] (
	.clk(CLK),
	.d(\PR|pc_id~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[21] .is_wysiwyg = "true";
defparam \prif.pc_id[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N3
dffeas \prif.pc_id[20] (
	.clk(CLK),
	.d(\PR|pc_id~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[20] .is_wysiwyg = "true";
defparam \prif.pc_id[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N17
dffeas \prif.pc_id[19] (
	.clk(CLK),
	.d(\PR|pc_id~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[19] .is_wysiwyg = "true";
defparam \prif.pc_id[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N15
dffeas \prif.pc_id[18] (
	.clk(CLK),
	.d(\PR|pc_id~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[18] .is_wysiwyg = "true";
defparam \prif.pc_id[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N1
dffeas \prif.pc_id[17] (
	.clk(CLK),
	.d(\PR|pc_id~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[17] .is_wysiwyg = "true";
defparam \prif.pc_id[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N23
dffeas \prif.pc_id[16] (
	.clk(CLK),
	.d(\PR|pc_id~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[16] .is_wysiwyg = "true";
defparam \prif.pc_id[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N13
dffeas \prif.pc_id[29] (
	.clk(CLK),
	.d(\PR|pc_id~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[29] .is_wysiwyg = "true";
defparam \prif.pc_id[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N19
dffeas \prif.pc_id[28] (
	.clk(CLK),
	.d(\PR|pc_id~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[28] .is_wysiwyg = "true";
defparam \prif.pc_id[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N1
dffeas \prif.pc_id[27] (
	.clk(CLK),
	.d(\PR|pc_id~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[27] .is_wysiwyg = "true";
defparam \prif.pc_id[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y32_N25
dffeas \prif.pc_id[26] (
	.clk(CLK),
	.d(\PR|pc_id~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[26] .is_wysiwyg = "true";
defparam \prif.pc_id[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y34_N27
dffeas \prif.pc_id[25] (
	.clk(CLK),
	.d(\PR|pc_id~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[25] .is_wysiwyg = "true";
defparam \prif.pc_id[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N15
dffeas \prif.pc_id[24] (
	.clk(CLK),
	.d(\PR|pc_id~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[24] .is_wysiwyg = "true";
defparam \prif.pc_id[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y34_N7
dffeas \prif.pc_id[31] (
	.clk(CLK),
	.d(\PR|pc_id~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[31] .is_wysiwyg = "true";
defparam \prif.pc_id[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y30_N29
dffeas \prif.pc_id[30] (
	.clk(CLK),
	.d(\PR|pc_id~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\HU|always1~5_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_id [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_id[30] .is_wysiwyg = "true";
defparam \prif.pc_id[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N4
cycloneive_lcell_comb \Add2~0 (
// Equation(s):
// \Add2~0_combout  = (pc_3 & (pc_2 $ (VCC))) # (!pc_3 & (pc_2 & VCC))
// \Add2~1  = CARRY((pc_3 & pc_2))

	.dataa(pc_3),
	.datab(pc_2),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add2~0_combout ),
	.cout(\Add2~1 ));
// synopsys translate_off
defparam \Add2~0 .lut_mask = 16'h6688;
defparam \Add2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N6
cycloneive_lcell_comb \Add2~2 (
// Equation(s):
// \Add2~2_combout  = (pc_4 & (!\Add2~1 )) # (!pc_4 & ((\Add2~1 ) # (GND)))
// \Add2~3  = CARRY((!\Add2~1 ) # (!pc_4))

	.dataa(gnd),
	.datab(pc_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~1 ),
	.combout(\Add2~2_combout ),
	.cout(\Add2~3 ));
// synopsys translate_off
defparam \Add2~2 .lut_mask = 16'h3C3F;
defparam \Add2~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N8
cycloneive_lcell_comb \Add2~4 (
// Equation(s):
// \Add2~4_combout  = (pc_5 & (\Add2~3  $ (GND))) # (!pc_5 & (!\Add2~3  & VCC))
// \Add2~5  = CARRY((pc_5 & !\Add2~3 ))

	.dataa(gnd),
	.datab(pc_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~3 ),
	.combout(\Add2~4_combout ),
	.cout(\Add2~5 ));
// synopsys translate_off
defparam \Add2~4 .lut_mask = 16'hC30C;
defparam \Add2~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N10
cycloneive_lcell_comb \Add2~6 (
// Equation(s):
// \Add2~6_combout  = (pc_6 & (!\Add2~5 )) # (!pc_6 & ((\Add2~5 ) # (GND)))
// \Add2~7  = CARRY((!\Add2~5 ) # (!pc_6))

	.dataa(gnd),
	.datab(pc_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~5 ),
	.combout(\Add2~6_combout ),
	.cout(\Add2~7 ));
// synopsys translate_off
defparam \Add2~6 .lut_mask = 16'h3C3F;
defparam \Add2~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N12
cycloneive_lcell_comb \Add2~8 (
// Equation(s):
// \Add2~8_combout  = (pc_7 & (\Add2~7  $ (GND))) # (!pc_7 & (!\Add2~7  & VCC))
// \Add2~9  = CARRY((pc_7 & !\Add2~7 ))

	.dataa(gnd),
	.datab(pc_7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~7 ),
	.combout(\Add2~8_combout ),
	.cout(\Add2~9 ));
// synopsys translate_off
defparam \Add2~8 .lut_mask = 16'hC30C;
defparam \Add2~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N14
cycloneive_lcell_comb \Add2~10 (
// Equation(s):
// \Add2~10_combout  = (pc_8 & (!\Add2~9 )) # (!pc_8 & ((\Add2~9 ) # (GND)))
// \Add2~11  = CARRY((!\Add2~9 ) # (!pc_8))

	.dataa(pc_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~9 ),
	.combout(\Add2~10_combout ),
	.cout(\Add2~11 ));
// synopsys translate_off
defparam \Add2~10 .lut_mask = 16'h5A5F;
defparam \Add2~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N16
cycloneive_lcell_comb \Add2~12 (
// Equation(s):
// \Add2~12_combout  = (pc_9 & (\Add2~11  $ (GND))) # (!pc_9 & (!\Add2~11  & VCC))
// \Add2~13  = CARRY((pc_9 & !\Add2~11 ))

	.dataa(pc_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~11 ),
	.combout(\Add2~12_combout ),
	.cout(\Add2~13 ));
// synopsys translate_off
defparam \Add2~12 .lut_mask = 16'hA50A;
defparam \Add2~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N18
cycloneive_lcell_comb \Add2~14 (
// Equation(s):
// \Add2~14_combout  = (pc_10 & (!\Add2~13 )) # (!pc_10 & ((\Add2~13 ) # (GND)))
// \Add2~15  = CARRY((!\Add2~13 ) # (!pc_10))

	.dataa(gnd),
	.datab(pc_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~13 ),
	.combout(\Add2~14_combout ),
	.cout(\Add2~15 ));
// synopsys translate_off
defparam \Add2~14 .lut_mask = 16'h3C3F;
defparam \Add2~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N20
cycloneive_lcell_comb \Add2~16 (
// Equation(s):
// \Add2~16_combout  = (pc_11 & (\Add2~15  $ (GND))) # (!pc_11 & (!\Add2~15  & VCC))
// \Add2~17  = CARRY((pc_11 & !\Add2~15 ))

	.dataa(gnd),
	.datab(pc_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~15 ),
	.combout(\Add2~16_combout ),
	.cout(\Add2~17 ));
// synopsys translate_off
defparam \Add2~16 .lut_mask = 16'hC30C;
defparam \Add2~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N22
cycloneive_lcell_comb \Add2~18 (
// Equation(s):
// \Add2~18_combout  = (pc_12 & (!\Add2~17 )) # (!pc_12 & ((\Add2~17 ) # (GND)))
// \Add2~19  = CARRY((!\Add2~17 ) # (!pc_12))

	.dataa(gnd),
	.datab(pc_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~17 ),
	.combout(\Add2~18_combout ),
	.cout(\Add2~19 ));
// synopsys translate_off
defparam \Add2~18 .lut_mask = 16'h3C3F;
defparam \Add2~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N24
cycloneive_lcell_comb \Add2~20 (
// Equation(s):
// \Add2~20_combout  = (pc_13 & (\Add2~19  $ (GND))) # (!pc_13 & (!\Add2~19  & VCC))
// \Add2~21  = CARRY((pc_13 & !\Add2~19 ))

	.dataa(pc_13),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~19 ),
	.combout(\Add2~20_combout ),
	.cout(\Add2~21 ));
// synopsys translate_off
defparam \Add2~20 .lut_mask = 16'hA50A;
defparam \Add2~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N26
cycloneive_lcell_comb \Add2~22 (
// Equation(s):
// \Add2~22_combout  = (pc_14 & (!\Add2~21 )) # (!pc_14 & ((\Add2~21 ) # (GND)))
// \Add2~23  = CARRY((!\Add2~21 ) # (!pc_14))

	.dataa(pc_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~21 ),
	.combout(\Add2~22_combout ),
	.cout(\Add2~23 ));
// synopsys translate_off
defparam \Add2~22 .lut_mask = 16'h5A5F;
defparam \Add2~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N28
cycloneive_lcell_comb \Add2~24 (
// Equation(s):
// \Add2~24_combout  = (pc_15 & (\Add2~23  $ (GND))) # (!pc_15 & (!\Add2~23  & VCC))
// \Add2~25  = CARRY((pc_15 & !\Add2~23 ))

	.dataa(gnd),
	.datab(pc_15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~23 ),
	.combout(\Add2~24_combout ),
	.cout(\Add2~25 ));
// synopsys translate_off
defparam \Add2~24 .lut_mask = 16'hC30C;
defparam \Add2~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N30
cycloneive_lcell_comb \Add2~26 (
// Equation(s):
// \Add2~26_combout  = (pc_16 & (!\Add2~25 )) # (!pc_16 & ((\Add2~25 ) # (GND)))
// \Add2~27  = CARRY((!\Add2~25 ) # (!pc_16))

	.dataa(pc_16),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~25 ),
	.combout(\Add2~26_combout ),
	.cout(\Add2~27 ));
// synopsys translate_off
defparam \Add2~26 .lut_mask = 16'h5A5F;
defparam \Add2~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N0
cycloneive_lcell_comb \Add2~28 (
// Equation(s):
// \Add2~28_combout  = (pc_17 & (\Add2~27  $ (GND))) # (!pc_17 & (!\Add2~27  & VCC))
// \Add2~29  = CARRY((pc_17 & !\Add2~27 ))

	.dataa(gnd),
	.datab(pc_17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~27 ),
	.combout(\Add2~28_combout ),
	.cout(\Add2~29 ));
// synopsys translate_off
defparam \Add2~28 .lut_mask = 16'hC30C;
defparam \Add2~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N2
cycloneive_lcell_comb \Add2~30 (
// Equation(s):
// \Add2~30_combout  = (pc_18 & (!\Add2~29 )) # (!pc_18 & ((\Add2~29 ) # (GND)))
// \Add2~31  = CARRY((!\Add2~29 ) # (!pc_18))

	.dataa(gnd),
	.datab(pc_18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~29 ),
	.combout(\Add2~30_combout ),
	.cout(\Add2~31 ));
// synopsys translate_off
defparam \Add2~30 .lut_mask = 16'h3C3F;
defparam \Add2~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N4
cycloneive_lcell_comb \Add2~32 (
// Equation(s):
// \Add2~32_combout  = (pc_19 & (\Add2~31  $ (GND))) # (!pc_19 & (!\Add2~31  & VCC))
// \Add2~33  = CARRY((pc_19 & !\Add2~31 ))

	.dataa(gnd),
	.datab(pc_19),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~31 ),
	.combout(\Add2~32_combout ),
	.cout(\Add2~33 ));
// synopsys translate_off
defparam \Add2~32 .lut_mask = 16'hC30C;
defparam \Add2~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N6
cycloneive_lcell_comb \Add2~34 (
// Equation(s):
// \Add2~34_combout  = (pc_20 & (!\Add2~33 )) # (!pc_20 & ((\Add2~33 ) # (GND)))
// \Add2~35  = CARRY((!\Add2~33 ) # (!pc_20))

	.dataa(gnd),
	.datab(pc_20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~33 ),
	.combout(\Add2~34_combout ),
	.cout(\Add2~35 ));
// synopsys translate_off
defparam \Add2~34 .lut_mask = 16'h3C3F;
defparam \Add2~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N8
cycloneive_lcell_comb \Add2~36 (
// Equation(s):
// \Add2~36_combout  = (pc_21 & (\Add2~35  $ (GND))) # (!pc_21 & (!\Add2~35  & VCC))
// \Add2~37  = CARRY((pc_21 & !\Add2~35 ))

	.dataa(pc_21),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~35 ),
	.combout(\Add2~36_combout ),
	.cout(\Add2~37 ));
// synopsys translate_off
defparam \Add2~36 .lut_mask = 16'hA50A;
defparam \Add2~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N10
cycloneive_lcell_comb \Add2~38 (
// Equation(s):
// \Add2~38_combout  = (pc_22 & (!\Add2~37 )) # (!pc_22 & ((\Add2~37 ) # (GND)))
// \Add2~39  = CARRY((!\Add2~37 ) # (!pc_22))

	.dataa(pc_22),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~37 ),
	.combout(\Add2~38_combout ),
	.cout(\Add2~39 ));
// synopsys translate_off
defparam \Add2~38 .lut_mask = 16'h5A5F;
defparam \Add2~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N12
cycloneive_lcell_comb \Add2~40 (
// Equation(s):
// \Add2~40_combout  = (pc_23 & (\Add2~39  $ (GND))) # (!pc_23 & (!\Add2~39  & VCC))
// \Add2~41  = CARRY((pc_23 & !\Add2~39 ))

	.dataa(pc_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~39 ),
	.combout(\Add2~40_combout ),
	.cout(\Add2~41 ));
// synopsys translate_off
defparam \Add2~40 .lut_mask = 16'hA50A;
defparam \Add2~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N14
cycloneive_lcell_comb \Add2~42 (
// Equation(s):
// \Add2~42_combout  = (pc_24 & (!\Add2~41 )) # (!pc_24 & ((\Add2~41 ) # (GND)))
// \Add2~43  = CARRY((!\Add2~41 ) # (!pc_24))

	.dataa(pc_24),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~41 ),
	.combout(\Add2~42_combout ),
	.cout(\Add2~43 ));
// synopsys translate_off
defparam \Add2~42 .lut_mask = 16'h5A5F;
defparam \Add2~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N16
cycloneive_lcell_comb \Add2~44 (
// Equation(s):
// \Add2~44_combout  = (pc_25 & (\Add2~43  $ (GND))) # (!pc_25 & (!\Add2~43  & VCC))
// \Add2~45  = CARRY((pc_25 & !\Add2~43 ))

	.dataa(gnd),
	.datab(pc_25),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~43 ),
	.combout(\Add2~44_combout ),
	.cout(\Add2~45 ));
// synopsys translate_off
defparam \Add2~44 .lut_mask = 16'hC30C;
defparam \Add2~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N18
cycloneive_lcell_comb \Add2~46 (
// Equation(s):
// \Add2~46_combout  = (pc_26 & (!\Add2~45 )) # (!pc_26 & ((\Add2~45 ) # (GND)))
// \Add2~47  = CARRY((!\Add2~45 ) # (!pc_26))

	.dataa(pc_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~45 ),
	.combout(\Add2~46_combout ),
	.cout(\Add2~47 ));
// synopsys translate_off
defparam \Add2~46 .lut_mask = 16'h5A5F;
defparam \Add2~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N20
cycloneive_lcell_comb \Add2~48 (
// Equation(s):
// \Add2~48_combout  = (pc_27 & (\Add2~47  $ (GND))) # (!pc_27 & (!\Add2~47  & VCC))
// \Add2~49  = CARRY((pc_27 & !\Add2~47 ))

	.dataa(gnd),
	.datab(pc_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~47 ),
	.combout(\Add2~48_combout ),
	.cout(\Add2~49 ));
// synopsys translate_off
defparam \Add2~48 .lut_mask = 16'hC30C;
defparam \Add2~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N22
cycloneive_lcell_comb \Add2~50 (
// Equation(s):
// \Add2~50_combout  = (pc_28 & (!\Add2~49 )) # (!pc_28 & ((\Add2~49 ) # (GND)))
// \Add2~51  = CARRY((!\Add2~49 ) # (!pc_28))

	.dataa(pc_28),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~49 ),
	.combout(\Add2~50_combout ),
	.cout(\Add2~51 ));
// synopsys translate_off
defparam \Add2~50 .lut_mask = 16'h5A5F;
defparam \Add2~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N24
cycloneive_lcell_comb \Add2~52 (
// Equation(s):
// \Add2~52_combout  = (pc_29 & (\Add2~51  $ (GND))) # (!pc_29 & (!\Add2~51  & VCC))
// \Add2~53  = CARRY((pc_29 & !\Add2~51 ))

	.dataa(gnd),
	.datab(pc_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~51 ),
	.combout(\Add2~52_combout ),
	.cout(\Add2~53 ));
// synopsys translate_off
defparam \Add2~52 .lut_mask = 16'hC30C;
defparam \Add2~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N26
cycloneive_lcell_comb \Add2~54 (
// Equation(s):
// \Add2~54_combout  = (pc_30 & (!\Add2~53 )) # (!pc_30 & ((\Add2~53 ) # (GND)))
// \Add2~55  = CARRY((!\Add2~53 ) # (!pc_30))

	.dataa(pc_30),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add2~53 ),
	.combout(\Add2~54_combout ),
	.cout(\Add2~55 ));
// synopsys translate_off
defparam \Add2~54 .lut_mask = 16'h5A5F;
defparam \Add2~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N28
cycloneive_lcell_comb \Add2~56 (
// Equation(s):
// \Add2~56_combout  = \Add2~55  $ (!pc_31)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(pc_31),
	.cin(\Add2~55 ),
	.combout(\Add2~56_combout ),
	.cout());
// synopsys translate_off
defparam \Add2~56 .lut_mask = 16'hF00F;
defparam \Add2~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X54_Y32_N15
dffeas \prif.ALUOP_ex[3] (
	.clk(CLK),
	.d(\PR|ALUOP_ex~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.ALUOP_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.ALUOP_ex[3] .is_wysiwyg = "true";
defparam \prif.ALUOP_ex[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N16
cycloneive_lcell_comb \Mux94~0 (
// Equation(s):
// \Mux94~0_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [1])))) # (!\prif.ALUScr_ex [0] & (\prif.shamt_ex [1] & ((\prif.ALUScr_ex [1]))))

	.dataa(\prif.shamt_ex [1]),
	.datab(\prif.imm_ex [1]),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\prif.ALUScr_ex [0]),
	.cin(gnd),
	.combout(\Mux94~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux94~0 .lut_mask = 16'hCCA0;
defparam \Mux94~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N30
cycloneive_lcell_comb \Mux89~2 (
// Equation(s):
// \Mux89~2_combout  = (!\prif.ALUScr_ex [1] & !\prif.ALUScr_ex [0])

	.dataa(gnd),
	.datab(gnd),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\prif.ALUScr_ex [0]),
	.cin(gnd),
	.combout(\Mux89~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux89~2 .lut_mask = 16'h000F;
defparam \Mux89~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y27_N3
dffeas \prif.Regwen_wb (
	.clk(CLK),
	.d(\PR|Regwen_wb~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.Regwen_wb~q ),
	.prn(vcc));
// synopsys translate_off
defparam \prif.Regwen_wb .is_wysiwyg = "true";
defparam \prif.Regwen_wb .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N29
dffeas \prif.regwrite_wb[2] (
	.clk(CLK),
	.d(\PR|regwrite_wb~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_wb [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_wb[2] .is_wysiwyg = "true";
defparam \prif.regwrite_wb[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N19
dffeas \prif.regwrite_wb[0] (
	.clk(CLK),
	.d(\PR|regwrite_wb~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_wb [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_wb[0] .is_wysiwyg = "true";
defparam \prif.regwrite_wb[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y27_N29
dffeas \prif.regwrite_wb[1] (
	.clk(CLK),
	.d(\PR|regwrite_wb~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_wb [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_wb[1] .is_wysiwyg = "true";
defparam \prif.regwrite_wb[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N25
dffeas \prif.regwrite_wb[4] (
	.clk(CLK),
	.d(\PR|regwrite_wb~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_wb [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_wb[4] .is_wysiwyg = "true";
defparam \prif.regwrite_wb[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y27_N15
dffeas \prif.regwrite_wb[3] (
	.clk(CLK),
	.d(\PR|regwrite_wb~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.regwrite_wb [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.regwrite_wb[3] .is_wysiwyg = "true";
defparam \prif.regwrite_wb[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N18
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (ptBScr & (prifdmemaddr_1 & !always01))

	.dataa(gnd),
	.datab(\HU|ptBScr~1_combout ),
	.datac(prifdmemaddr_1),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'h00C0;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y28_N23
dffeas \prif.dmemload_wb[1] (
	.clk(CLK),
	.d(\PR|dmemload_wb~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[1] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y28_N21
dffeas \prif.dmemaddr_wb[1] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[1] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N7
dffeas \prif.dataScr_wb[0] (
	.clk(CLK),
	.d(\PR|dataScr_wb~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dataScr_wb [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dataScr_wb[0] .is_wysiwyg = "true";
defparam \prif.dataScr_wb[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N29
dffeas \prif.dataScr_wb[1] (
	.clk(CLK),
	.d(\PR|dataScr_wb~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dataScr_wb [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dataScr_wb[1] .is_wysiwyg = "true";
defparam \prif.dataScr_wb[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N14
cycloneive_lcell_comb \Mux163~0 (
// Equation(s):
// \Mux163~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [1])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [1])))))

	.dataa(\prif.dmemload_wb [1]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dmemaddr_wb [1]),
	.cin(gnd),
	.combout(\Mux163~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux163~0 .lut_mask = 16'h0B08;
defparam \Mux163~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y28_N3
dffeas \prif.pc_wb[1] (
	.clk(CLK),
	.d(\PR|pc_wb~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[1] .is_wysiwyg = "true";
defparam \prif.pc_wb[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N8
cycloneive_lcell_comb \Mux163~1 (
// Equation(s):
// \Mux163~1_combout  = (\Mux163~0_combout ) # ((\prif.dataScr_wb [1] & (\prif.dataScr_wb [0] & \prif.pc_wb [1])))

	.dataa(\Mux163~0_combout ),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dataScr_wb [0]),
	.datad(\prif.pc_wb [1]),
	.cin(gnd),
	.combout(\Mux163~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux163~1 .lut_mask = 16'hEAAA;
defparam \Mux163~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N14
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (!ptBScr & ((always01 & ((\Mux163~1_combout ))) # (!always01 & (\prif.rdat2_ex [1]))))

	.dataa(\HU|always0~5_combout ),
	.datab(\prif.rdat2_ex [1]),
	.datac(\Mux163~1_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'h00E4;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N12
cycloneive_lcell_comb \Mux94~1 (
// Equation(s):
// \Mux94~1_combout  = (\Mux94~0_combout ) # ((\Mux89~2_combout  & ((\Mux62~1_combout ) # (\Mux62~0_combout ))))

	.dataa(\Mux62~1_combout ),
	.datab(\Mux94~0_combout ),
	.datac(\Mux89~2_combout ),
	.datad(\Mux62~0_combout ),
	.cin(gnd),
	.combout(\Mux94~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux94~1 .lut_mask = 16'hFCEC;
defparam \Mux94~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y27_N27
dffeas \prif.rs_ex[1] (
	.clk(CLK),
	.d(\PR|prif.rs_ex[1]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rs_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rs_ex[1] .is_wysiwyg = "true";
defparam \prif.rs_ex[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y27_N17
dffeas \prif.rs_ex[0] (
	.clk(CLK),
	.d(\PR|prif.rs_ex[0]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rs_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rs_ex[0] .is_wysiwyg = "true";
defparam \prif.rs_ex[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y27_N21
dffeas \prif.rs_ex[3] (
	.clk(CLK),
	.d(\PR|prif.rs_ex[3]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rs_ex [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rs_ex[3] .is_wysiwyg = "true";
defparam \prif.rs_ex[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y27_N31
dffeas \prif.rs_ex[2] (
	.clk(CLK),
	.d(\PR|prif.rs_ex[2]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rs_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rs_ex[2] .is_wysiwyg = "true";
defparam \prif.rs_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y27_N7
dffeas \prif.rs_ex[4] (
	.clk(CLK),
	.d(\PR|prif.rs_ex[4]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rs_ex [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rs_ex[4] .is_wysiwyg = "true";
defparam \prif.rs_ex[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N12
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (always02 & ((prifdmemaddr_1))) # (!always02 & (\prif.rdat1_ex [1]))

	.dataa(gnd),
	.datab(\prif.rdat1_ex [1]),
	.datac(prifdmemaddr_1),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hF0CC;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N22
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (ptAScr & (((\Mux163~1_combout  & !always02)))) # (!ptAScr & (\Mux30~0_combout ))

	.dataa(\Mux30~0_combout ),
	.datab(\Mux163~1_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'h0CAA;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N20
cycloneive_lcell_comb \Mux95~0 (
// Equation(s):
// \Mux95~0_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [0])))) # (!\prif.ALUScr_ex [0] & (\prif.shamt_ex [0] & (\prif.ALUScr_ex [1])))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.shamt_ex [0]),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\prif.imm_ex [0]),
	.cin(gnd),
	.combout(\Mux95~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux95~0 .lut_mask = 16'hEA40;
defparam \Mux95~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N6
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (!always01 & (prifdmemaddr_0 & ptBScr))

	.dataa(gnd),
	.datab(\HU|always0~5_combout ),
	.datac(prifdmemaddr_0),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'h3000;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y28_N19
dffeas \prif.dmemload_wb[0] (
	.clk(CLK),
	.d(\PR|dmemload_wb~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[0] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y28_N21
dffeas \prif.dmemaddr_wb[0] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[0] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N6
cycloneive_lcell_comb \Mux164~0 (
// Equation(s):
// \Mux164~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [0]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [0]))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dmemaddr_wb [0]),
	.datac(\prif.dataScr_wb [0]),
	.datad(\prif.dmemload_wb [0]),
	.cin(gnd),
	.combout(\Mux164~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux164~0 .lut_mask = 16'h5404;
defparam \Mux164~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y28_N1
dffeas \prif.pc_wb[0] (
	.clk(CLK),
	.d(\PR|pc_wb~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[0] .is_wysiwyg = "true";
defparam \prif.pc_wb[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N22
cycloneive_lcell_comb \Mux164~1 (
// Equation(s):
// \Mux164~1_combout  = (\Mux164~0_combout ) # ((\prif.dataScr_wb [1] & (\prif.dataScr_wb [0] & \prif.pc_wb [0])))

	.dataa(\Mux164~0_combout ),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dataScr_wb [0]),
	.datad(\prif.pc_wb [0]),
	.cin(gnd),
	.combout(\Mux164~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux164~1 .lut_mask = 16'hEAAA;
defparam \Mux164~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N8
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (!ptBScr & ((always01 & (\Mux164~1_combout )) # (!always01 & ((\prif.rdat2_ex [0])))))

	.dataa(\Mux164~1_combout ),
	.datab(\prif.rdat2_ex [0]),
	.datac(\HU|always0~5_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'h00AC;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N26
cycloneive_lcell_comb \Mux95~1 (
// Equation(s):
// \Mux95~1_combout  = (\Mux95~0_combout ) # ((\Mux89~2_combout  & ((\Mux63~1_combout ) # (\Mux63~0_combout ))))

	.dataa(\Mux89~2_combout ),
	.datab(\Mux95~0_combout ),
	.datac(\Mux63~1_combout ),
	.datad(\Mux63~0_combout ),
	.cin(gnd),
	.combout(\Mux95~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux95~1 .lut_mask = 16'hEEEC;
defparam \Mux95~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N0
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (always02 & ((prifdmemaddr_0))) # (!always02 & (\prif.rdat1_ex [0]))

	.dataa(\prif.rdat1_ex [0]),
	.datab(gnd),
	.datac(prifdmemaddr_0),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hF0AA;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N14
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (ptAScr & (!always02 & (\Mux164~1_combout ))) # (!ptAScr & (((\Mux31~0_combout ))))

	.dataa(\HU|always0~6_combout ),
	.datab(\HU|ptAScr~4_combout ),
	.datac(\Mux164~1_combout ),
	.datad(\Mux31~0_combout ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'h7340;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y27_N13
dffeas \prif.dmemload_wb[3] (
	.clk(CLK),
	.d(\PR|dmemload_wb~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[3] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y27_N27
dffeas \prif.dmemaddr_wb[3] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[3] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N4
cycloneive_lcell_comb \Mux161~0 (
// Equation(s):
// \Mux161~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [3]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [3]))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.dmemaddr_wb [3]),
	.datad(\prif.dmemload_wb [3]),
	.cin(gnd),
	.combout(\Mux161~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux161~0 .lut_mask = 16'h5410;
defparam \Mux161~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y27_N11
dffeas \prif.pc_wb[3] (
	.clk(CLK),
	.d(\PR|pc_wb~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[3] .is_wysiwyg = "true";
defparam \prif.pc_wb[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N20
cycloneive_lcell_comb \Mux161~1 (
// Equation(s):
// \Mux161~1_combout  = (\Mux161~0_combout ) # ((\prif.dataScr_wb [1] & (\prif.dataScr_wb [0] & \prif.pc_wb [3])))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\Mux161~0_combout ),
	.datad(\prif.pc_wb [3]),
	.cin(gnd),
	.combout(\Mux161~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux161~1 .lut_mask = 16'hF8F0;
defparam \Mux161~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N12
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (!ptBScr & ((always01 & (\Mux161~1_combout )) # (!always01 & ((\prif.rdat2_ex [3])))))

	.dataa(\Mux161~1_combout ),
	.datab(\prif.rdat2_ex [3]),
	.datac(\HU|always0~5_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'h00AC;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N22
cycloneive_lcell_comb \Mux92~0 (
// Equation(s):
// \Mux92~0_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [3])))) # (!\prif.ALUScr_ex [0] & (\prif.shamt_ex [3] & (\prif.ALUScr_ex [1])))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.shamt_ex [3]),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\prif.imm_ex [3]),
	.cin(gnd),
	.combout(\Mux92~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux92~0 .lut_mask = 16'hEA40;
defparam \Mux92~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N24
cycloneive_lcell_comb \Mux92~1 (
// Equation(s):
// \Mux92~1_combout  = (!always01 & (prifdmemaddr_3 & ptBScr))

	.dataa(gnd),
	.datab(\HU|always0~5_combout ),
	.datac(prifdmemaddr_3),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux92~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux92~1 .lut_mask = 16'h3000;
defparam \Mux92~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N14
cycloneive_lcell_comb \Mux92~2 (
// Equation(s):
// \Mux92~2_combout  = (\Mux92~0_combout ) # ((\Mux89~2_combout  & ((\Mux92~1_combout ) # (\Mux60~0_combout ))))

	.dataa(\Mux92~0_combout ),
	.datab(\Mux92~1_combout ),
	.datac(\Mux89~2_combout ),
	.datad(\Mux60~0_combout ),
	.cin(gnd),
	.combout(\Mux92~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux92~2 .lut_mask = 16'hFAEA;
defparam \Mux92~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N22
cycloneive_lcell_comb \Mux93~0 (
// Equation(s):
// \Mux93~0_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [2])))) # (!\prif.ALUScr_ex [0] & (\prif.ALUScr_ex [1] & (\prif.shamt_ex [2])))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.shamt_ex [2]),
	.datac(\prif.imm_ex [2]),
	.datad(\prif.ALUScr_ex [0]),
	.cin(gnd),
	.combout(\Mux93~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux93~0 .lut_mask = 16'hF088;
defparam \Mux93~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y29_N7
dffeas \prif.dmemload_wb[2] (
	.clk(CLK),
	.d(\PR|dmemload_wb~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[2] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y29_N5
dffeas \prif.dmemaddr_wb[2] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[2] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N30
cycloneive_lcell_comb \Mux162~0 (
// Equation(s):
// \Mux162~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [2]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [2]))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dmemaddr_wb [2]),
	.datad(\prif.dmemload_wb [2]),
	.cin(gnd),
	.combout(\Mux162~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux162~0 .lut_mask = 16'h3210;
defparam \Mux162~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y29_N29
dffeas \prif.pc_wb[2] (
	.clk(CLK),
	.d(\PR|pc_wb~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[2] .is_wysiwyg = "true";
defparam \prif.pc_wb[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N14
cycloneive_lcell_comb \Mux162~1 (
// Equation(s):
// \Mux162~1_combout  = (\Mux162~0_combout ) # ((\prif.dataScr_wb [0] & (\prif.dataScr_wb [1] & \prif.pc_wb [2])))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\Mux162~0_combout ),
	.datad(\prif.pc_wb [2]),
	.cin(gnd),
	.combout(\Mux162~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux162~1 .lut_mask = 16'hF8F0;
defparam \Mux162~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N24
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (!ptBScr & ((always01 & (\Mux162~1_combout )) # (!always01 & ((\prif.rdat2_ex [2])))))

	.dataa(\Mux162~1_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(\prif.rdat2_ex [2]),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'h00B8;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N26
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (\Mux61~0_combout ) # ((ptBScr & (prifdmemaddr_2 & !always01)))

	.dataa(\Mux61~0_combout ),
	.datab(\HU|ptBScr~1_combout ),
	.datac(prifdmemaddr_2),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hAAEA;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y27_N23
dffeas \prif.dmemload_wb[4] (
	.clk(CLK),
	.d(\PR|dmemload_wb~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[4] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y27_N17
dffeas \prif.dmemaddr_wb[4] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[4] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N18
cycloneive_lcell_comb \Mux160~0 (
// Equation(s):
// \Mux160~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [4])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [4])))))

	.dataa(\prif.dmemload_wb [4]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dmemaddr_wb [4]),
	.cin(gnd),
	.combout(\Mux160~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux160~0 .lut_mask = 16'h0B08;
defparam \Mux160~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y27_N9
dffeas \prif.pc_wb[4] (
	.clk(CLK),
	.d(\PR|pc_wb~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[4] .is_wysiwyg = "true";
defparam \prif.pc_wb[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N30
cycloneive_lcell_comb \Mux160~1 (
// Equation(s):
// \Mux160~1_combout  = (\Mux160~0_combout ) # ((\prif.dataScr_wb [1] & (\prif.dataScr_wb [0] & \prif.pc_wb [4])))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.pc_wb [4]),
	.datad(\Mux160~0_combout ),
	.cin(gnd),
	.combout(\Mux160~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux160~1 .lut_mask = 16'hFF80;
defparam \Mux160~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N24
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (!ptBScr & ((always01 & ((\Mux160~1_combout ))) # (!always01 & (\prif.rdat2_ex [4]))))

	.dataa(\prif.rdat2_ex [4]),
	.datab(\HU|always0~5_combout ),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\Mux160~1_combout ),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'h0E02;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N18
cycloneive_lcell_comb \Mux91~0 (
// Equation(s):
// \Mux91~0_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [4])))) # (!\prif.ALUScr_ex [0] & (\prif.ALUScr_ex [1] & (\prif.shamt_ex [4])))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.ALUScr_ex [1]),
	.datac(\prif.shamt_ex [4]),
	.datad(\prif.imm_ex [4]),
	.cin(gnd),
	.combout(\Mux91~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux91~0 .lut_mask = 16'hEA40;
defparam \Mux91~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N26
cycloneive_lcell_comb \Mux91~1 (
// Equation(s):
// \Mux91~1_combout  = (ptBScr & (!always01 & prifdmemaddr_4))

	.dataa(gnd),
	.datab(\HU|ptBScr~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(prifdmemaddr_4),
	.cin(gnd),
	.combout(\Mux91~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux91~1 .lut_mask = 16'h0C00;
defparam \Mux91~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N20
cycloneive_lcell_comb \Mux91~2 (
// Equation(s):
// \Mux91~2_combout  = (\Mux91~0_combout ) # ((\Mux89~2_combout  & ((\Mux59~0_combout ) # (\Mux91~1_combout ))))

	.dataa(\Mux89~2_combout ),
	.datab(\Mux59~0_combout ),
	.datac(\Mux91~1_combout ),
	.datad(\Mux91~0_combout ),
	.cin(gnd),
	.combout(\Mux91~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux91~2 .lut_mask = 16'hFFA8;
defparam \Mux91~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y28_N13
dffeas \prif.dmemload_wb[31] (
	.clk(CLK),
	.d(\PR|dmemload_wb~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[31] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N27
dffeas \prif.imm_wb[15] (
	.clk(CLK),
	.d(\PR|imm_wb~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[15] .is_wysiwyg = "true";
defparam \prif.imm_wb[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N17
dffeas \prif.dmemaddr_wb[31] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[31] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N6
cycloneive_lcell_comb \Mux133~0 (
// Equation(s):
// \Mux133~0_combout  = (\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0]) # ((\prif.imm_wb [15])))) # (!\prif.dataScr_wb [1] & (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [31]))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.imm_wb [15]),
	.datad(\prif.dmemaddr_wb [31]),
	.cin(gnd),
	.combout(\Mux133~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux133~0 .lut_mask = 16'hB9A8;
defparam \Mux133~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y28_N5
dffeas \prif.pc_wb[31] (
	.clk(CLK),
	.d(\PR|pc_wb~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[31] .is_wysiwyg = "true";
defparam \prif.pc_wb[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N10
cycloneive_lcell_comb \Mux133~1 (
// Equation(s):
// \Mux133~1_combout  = (\prif.dataScr_wb [0] & ((\Mux133~0_combout  & ((\prif.pc_wb [31]))) # (!\Mux133~0_combout  & (\prif.dmemload_wb [31])))) # (!\prif.dataScr_wb [0] & (((\Mux133~0_combout ))))

	.dataa(\prif.dmemload_wb [31]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.pc_wb [31]),
	.datad(\Mux133~0_combout ),
	.cin(gnd),
	.combout(\Mux133~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux133~1 .lut_mask = 16'hF388;
defparam \Mux133~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N14
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (ptBScr & (((prifdmemaddr_31) # (always01)))) # (!ptBScr & (\prif.rdat2_ex [31] & ((!always01))))

	.dataa(\prif.rdat2_ex [31]),
	.datab(prifdmemaddr_31),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hF0CA;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N24
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (\Mux32~0_combout  & ((\prif.imm_mem [15]) # ((!always01)))) # (!\Mux32~0_combout  & (((\Mux133~1_combout  & always01))))

	.dataa(\prif.imm_mem [15]),
	.datab(\Mux32~0_combout ),
	.datac(\Mux133~1_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hB8CC;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N30
cycloneive_lcell_comb \Mux64~0 (
// Equation(s):
// \Mux64~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux32~1_combout )))))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.instr_ex [15]),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\Mux32~1_combout ),
	.cin(gnd),
	.combout(\Mux64~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux64~0 .lut_mask = 16'h0D08;
defparam \Mux64~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y28_N17
dffeas \prif.imm_wb[14] (
	.clk(CLK),
	.d(\PR|imm_wb~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[14] .is_wysiwyg = "true";
defparam \prif.imm_wb[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N31
dffeas \prif.dmemload_wb[30] (
	.clk(CLK),
	.d(\PR|dmemload_wb~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[30] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N21
dffeas \prif.dmemaddr_wb[30] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[30] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N18
cycloneive_lcell_comb \Mux134~0 (
// Equation(s):
// \Mux134~0_combout  = (\prif.dataScr_wb [0] & ((\prif.dmemload_wb [30]) # ((\prif.dataScr_wb [1])))) # (!\prif.dataScr_wb [0] & (((\prif.dmemaddr_wb [30] & !\prif.dataScr_wb [1]))))

	.dataa(\prif.dmemload_wb [30]),
	.datab(\prif.dmemaddr_wb [30]),
	.datac(\prif.dataScr_wb [0]),
	.datad(\prif.dataScr_wb [1]),
	.cin(gnd),
	.combout(\Mux134~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux134~0 .lut_mask = 16'hF0AC;
defparam \Mux134~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y28_N5
dffeas \prif.pc_wb[30] (
	.clk(CLK),
	.d(\PR|pc_wb~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[30] .is_wysiwyg = "true";
defparam \prif.pc_wb[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N10
cycloneive_lcell_comb \Mux134~1 (
// Equation(s):
// \Mux134~1_combout  = (\prif.dataScr_wb [1] & ((\Mux134~0_combout  & (\prif.pc_wb [30])) # (!\Mux134~0_combout  & ((\prif.imm_wb [14]))))) # (!\prif.dataScr_wb [1] & (\Mux134~0_combout ))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\Mux134~0_combout ),
	.datac(\prif.pc_wb [30]),
	.datad(\prif.imm_wb [14]),
	.cin(gnd),
	.combout(\Mux134~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux134~1 .lut_mask = 16'hE6C4;
defparam \Mux134~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N8
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (always01 & ((\Mux134~1_combout ) # ((ptBScr)))) # (!always01 & (((\prif.rdat2_ex [30] & !ptBScr))))

	.dataa(\Mux134~1_combout ),
	.datab(\prif.rdat2_ex [30]),
	.datac(\HU|always0~5_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hF0AC;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N14
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (\Mux33~0_combout  & ((\prif.imm_mem [14]) # ((!ptBScr)))) # (!\Mux33~0_combout  & (((prifdmemaddr_30 & ptBScr))))

	.dataa(\prif.imm_mem [14]),
	.datab(prifdmemaddr_30),
	.datac(\Mux33~0_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hACF0;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N24
cycloneive_lcell_comb \Mux65~0 (
// Equation(s):
// \Mux65~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & ((\prif.instr_ex [15]))) # (!\prif.ALUScr_ex [0] & (\Mux33~1_combout ))))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.ALUScr_ex [1]),
	.datac(\Mux33~1_combout ),
	.datad(\prif.instr_ex [15]),
	.cin(gnd),
	.combout(\Mux65~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux65~0 .lut_mask = 16'h3210;
defparam \Mux65~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N23
dffeas \prif.dmemload_wb[29] (
	.clk(CLK),
	.d(\PR|dmemload_wb~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[29] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N13
dffeas \prif.imm_wb[13] (
	.clk(CLK),
	.d(\PR|imm_wb~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[13] .is_wysiwyg = "true";
defparam \prif.imm_wb[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N11
dffeas \prif.dmemaddr_wb[29] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[29] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N20
cycloneive_lcell_comb \Mux135~0 (
// Equation(s):
// \Mux135~0_combout  = (\prif.dataScr_wb [1] & (((\prif.dataScr_wb [0]) # (\prif.imm_wb [13])))) # (!\prif.dataScr_wb [1] & (\prif.dmemaddr_wb [29] & (!\prif.dataScr_wb [0])))

	.dataa(\prif.dmemaddr_wb [29]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dataScr_wb [0]),
	.datad(\prif.imm_wb [13]),
	.cin(gnd),
	.combout(\Mux135~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux135~0 .lut_mask = 16'hCEC2;
defparam \Mux135~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N15
dffeas \prif.pc_wb[29] (
	.clk(CLK),
	.d(\PR|pc_wb~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[29] .is_wysiwyg = "true";
defparam \prif.pc_wb[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N16
cycloneive_lcell_comb \Mux135~1 (
// Equation(s):
// \Mux135~1_combout  = (\prif.dataScr_wb [0] & ((\Mux135~0_combout  & ((\prif.pc_wb [29]))) # (!\Mux135~0_combout  & (\prif.dmemload_wb [29])))) # (!\prif.dataScr_wb [0] & (((\Mux135~0_combout ))))

	.dataa(\prif.dmemload_wb [29]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.pc_wb [29]),
	.datad(\Mux135~0_combout ),
	.cin(gnd),
	.combout(\Mux135~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux135~1 .lut_mask = 16'hF388;
defparam \Mux135~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N30
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (ptBScr & ((always01) # ((prifdmemaddr_29)))) # (!ptBScr & (!always01 & ((\prif.rdat2_ex [29]))))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(prifdmemaddr_29),
	.datad(\prif.rdat2_ex [29]),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hB9A8;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N28
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (always01 & ((\Mux34~0_combout  & ((\prif.imm_mem [13]))) # (!\Mux34~0_combout  & (\Mux135~1_combout )))) # (!always01 & (((\Mux34~0_combout ))))

	.dataa(\Mux135~1_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(\Mux34~0_combout ),
	.datad(\prif.imm_mem [13]),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hF838;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N2
cycloneive_lcell_comb \Mux66~0 (
// Equation(s):
// \Mux66~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux34~1_combout )))))

	.dataa(\prif.instr_ex [15]),
	.datab(\prif.ALUScr_ex [1]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux34~1_combout ),
	.cin(gnd),
	.combout(\Mux66~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux66~0 .lut_mask = 16'h2320;
defparam \Mux66~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y28_N21
dffeas \prif.dmemload_wb[5] (
	.clk(CLK),
	.d(\PR|dmemload_wb~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[5] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y28_N23
dffeas \prif.dmemaddr_wb[5] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[5] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N28
cycloneive_lcell_comb \Mux159~0 (
// Equation(s):
// \Mux159~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [5]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [5]))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.dmemaddr_wb [5]),
	.datad(\prif.dmemload_wb [5]),
	.cin(gnd),
	.combout(\Mux159~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux159~0 .lut_mask = 16'h5410;
defparam \Mux159~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y31_N13
dffeas \prif.pc_wb[5] (
	.clk(CLK),
	.d(\PR|pc_wb~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[5] .is_wysiwyg = "true";
defparam \prif.pc_wb[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N14
cycloneive_lcell_comb \Mux159~1 (
// Equation(s):
// \Mux159~1_combout  = (\Mux159~0_combout ) # ((\prif.dataScr_wb [1] & (\prif.pc_wb [5] & \prif.dataScr_wb [0])))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\Mux159~0_combout ),
	.datac(\prif.pc_wb [5]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux159~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux159~1 .lut_mask = 16'hECCC;
defparam \Mux159~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N12
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (!ptBScr & ((always01 & (\Mux159~1_combout )) # (!always01 & ((\prif.rdat2_ex [5])))))

	.dataa(\Mux159~1_combout ),
	.datab(\prif.rdat2_ex [5]),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'h0A0C;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N2
cycloneive_lcell_comb \Mux90~2 (
// Equation(s):
// \Mux90~2_combout  = (\Mux58~0_combout ) # ((prifdmemaddr_5 & (ptBScr & !always01)))

	.dataa(\Mux58~0_combout ),
	.datab(prifdmemaddr_5),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux90~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux90~2 .lut_mask = 16'hAAEA;
defparam \Mux90~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y29_N31
dffeas \prif.dmemload_wb[15] (
	.clk(CLK),
	.d(\PR|dmemload_wb~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[15] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y26_N3
dffeas \prif.dmemaddr_wb[15] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[15] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N12
cycloneive_lcell_comb \Mux149~0 (
// Equation(s):
// \Mux149~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [15])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [15])))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dmemload_wb [15]),
	.datad(\prif.dmemaddr_wb [15]),
	.cin(gnd),
	.combout(\Mux149~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux149~0 .lut_mask = 16'h3120;
defparam \Mux149~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y29_N27
dffeas \prif.pc_wb[15] (
	.clk(CLK),
	.d(\PR|pc_wb~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[15] .is_wysiwyg = "true";
defparam \prif.pc_wb[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N16
cycloneive_lcell_comb \Mux149~1 (
// Equation(s):
// \Mux149~1_combout  = (\Mux149~0_combout ) # ((\prif.dataScr_wb [0] & (\prif.dataScr_wb [1] & \prif.pc_wb [15])))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.pc_wb [15]),
	.datad(\Mux149~0_combout ),
	.cin(gnd),
	.combout(\Mux149~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux149~1 .lut_mask = 16'hFF80;
defparam \Mux149~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N12
cycloneive_lcell_comb \Mux80~2 (
// Equation(s):
// \Mux80~2_combout  = (ptBScr & (((always01)))) # (!ptBScr & ((always01 & ((\Mux149~1_combout ))) # (!always01 & (\prif.rdat2_ex [15]))))

	.dataa(\prif.rdat2_ex [15]),
	.datab(\HU|ptBScr~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux149~1_combout ),
	.cin(gnd),
	.combout(\Mux80~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux80~2 .lut_mask = 16'hF2C2;
defparam \Mux80~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N18
cycloneive_lcell_comb \Mux80~3 (
// Equation(s):
// \Mux80~3_combout  = (\Mux80~2_combout  & ((!ptBScr))) # (!\Mux80~2_combout  & (prifdmemaddr_15 & ptBScr))

	.dataa(\Mux80~2_combout ),
	.datab(gnd),
	.datac(prifdmemaddr_15),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux80~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux80~3 .lut_mask = 16'h50AA;
defparam \Mux80~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y26_N23
dffeas \prif.dmemload_wb[14] (
	.clk(CLK),
	.d(\PR|dmemload_wb~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[14] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y26_N25
dffeas \prif.dmemaddr_wb[14] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[14] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N14
cycloneive_lcell_comb \Mux150~0 (
// Equation(s):
// \Mux150~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [14]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [14]))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dmemaddr_wb [14]),
	.datac(\prif.dmemload_wb [14]),
	.datad(\prif.dataScr_wb [1]),
	.cin(gnd),
	.combout(\Mux150~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux150~0 .lut_mask = 16'h00E4;
defparam \Mux150~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y26_N29
dffeas \prif.pc_wb[14] (
	.clk(CLK),
	.d(\PR|pc_wb~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[14] .is_wysiwyg = "true";
defparam \prif.pc_wb[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N26
cycloneive_lcell_comb \Mux150~1 (
// Equation(s):
// \Mux150~1_combout  = (\Mux150~0_combout ) # ((\prif.dataScr_wb [1] & (\prif.pc_wb [14] & \prif.dataScr_wb [0])))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.pc_wb [14]),
	.datac(\Mux150~0_combout ),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux150~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux150~1 .lut_mask = 16'hF8F0;
defparam \Mux150~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N12
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (!ptBScr & ((always01 & (\Mux150~1_combout )) # (!always01 & ((\prif.rdat2_ex [14])))))

	.dataa(\Mux150~1_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\prif.rdat2_ex [14]),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'h0B08;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N10
cycloneive_lcell_comb \Mux81~2 (
// Equation(s):
// \Mux81~2_combout  = (\Mux49~0_combout ) # ((ptBScr & (prifdmemaddr_14 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_14),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux49~0_combout ),
	.cin(gnd),
	.combout(\Mux81~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux81~2 .lut_mask = 16'hFF08;
defparam \Mux81~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y26_N13
dffeas \prif.dmemload_wb[13] (
	.clk(CLK),
	.d(\PR|dmemload_wb~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[13] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y26_N3
dffeas \prif.dmemaddr_wb[13] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[13] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N24
cycloneive_lcell_comb \Mux151~0 (
// Equation(s):
// \Mux151~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [13]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [13]))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dmemaddr_wb [13]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dmemload_wb [13]),
	.cin(gnd),
	.combout(\Mux151~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux151~0 .lut_mask = 16'h0E04;
defparam \Mux151~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y26_N23
dffeas \prif.pc_wb[13] (
	.clk(CLK),
	.d(\PR|pc_wb~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[13] .is_wysiwyg = "true";
defparam \prif.pc_wb[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N16
cycloneive_lcell_comb \Mux151~1 (
// Equation(s):
// \Mux151~1_combout  = (\Mux151~0_combout ) # ((\prif.dataScr_wb [1] & (\prif.pc_wb [13] & \prif.dataScr_wb [0])))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\Mux151~0_combout ),
	.datac(\prif.pc_wb [13]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux151~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux151~1 .lut_mask = 16'hECCC;
defparam \Mux151~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N10
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (!ptBScr & ((always01 & ((\Mux151~1_combout ))) # (!always01 & (\prif.rdat2_ex [13]))))

	.dataa(\prif.rdat2_ex [13]),
	.datab(\HU|ptBScr~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux151~1_combout ),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'h3202;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N0
cycloneive_lcell_comb \Mux82~2 (
// Equation(s):
// \Mux82~2_combout  = (\Mux50~0_combout ) # ((!always01 & (ptBScr & prifdmemaddr_13)))

	.dataa(\HU|always0~5_combout ),
	.datab(\HU|ptBScr~1_combout ),
	.datac(prifdmemaddr_13),
	.datad(\Mux50~0_combout ),
	.cin(gnd),
	.combout(\Mux82~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux82~2 .lut_mask = 16'hFF40;
defparam \Mux82~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y28_N21
dffeas \prif.dmemload_wb[12] (
	.clk(CLK),
	.d(\PR|dmemload_wb~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[12] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y28_N31
dffeas \prif.dmemaddr_wb[12] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[12] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N4
cycloneive_lcell_comb \Mux152~0 (
// Equation(s):
// \Mux152~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [12])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [12])))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dmemload_wb [12]),
	.datac(\prif.dmemaddr_wb [12]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux152~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux152~0 .lut_mask = 16'h4450;
defparam \Mux152~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y28_N27
dffeas \prif.pc_wb[12] (
	.clk(CLK),
	.d(\PR|pc_wb~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[12] .is_wysiwyg = "true";
defparam \prif.pc_wb[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N8
cycloneive_lcell_comb \Mux152~1 (
// Equation(s):
// \Mux152~1_combout  = (\Mux152~0_combout ) # ((\prif.pc_wb [12] & (\prif.dataScr_wb [0] & \prif.dataScr_wb [1])))

	.dataa(\prif.pc_wb [12]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\Mux152~0_combout ),
	.datad(\prif.dataScr_wb [1]),
	.cin(gnd),
	.combout(\Mux152~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux152~1 .lut_mask = 16'hF8F0;
defparam \Mux152~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N2
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (!ptBScr & ((always01 & ((\Mux152~1_combout ))) # (!always01 & (\prif.rdat2_ex [12]))))

	.dataa(\prif.rdat2_ex [12]),
	.datab(\HU|always0~5_combout ),
	.datac(\Mux152~1_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'h00E2;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N24
cycloneive_lcell_comb \Mux83~2 (
// Equation(s):
// \Mux83~2_combout  = (\Mux51~0_combout ) # ((ptBScr & (prifdmemaddr_12 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_12),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux51~0_combout ),
	.cin(gnd),
	.combout(\Mux83~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux83~2 .lut_mask = 16'hFF08;
defparam \Mux83~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y28_N7
dffeas \prif.dmemload_wb[11] (
	.clk(CLK),
	.d(\PR|dmemload_wb~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[11] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y28_N29
dffeas \prif.dmemaddr_wb[11] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[11] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N18
cycloneive_lcell_comb \Mux153~0 (
// Equation(s):
// \Mux153~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [11])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [11])))))

	.dataa(\prif.dmemload_wb [11]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dataScr_wb [0]),
	.datad(\prif.dmemaddr_wb [11]),
	.cin(gnd),
	.combout(\Mux153~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux153~0 .lut_mask = 16'h2320;
defparam \Mux153~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y28_N9
dffeas \prif.pc_wb[11] (
	.clk(CLK),
	.d(\PR|pc_wb~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[11] .is_wysiwyg = "true";
defparam \prif.pc_wb[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N2
cycloneive_lcell_comb \Mux153~1 (
// Equation(s):
// \Mux153~1_combout  = (\Mux153~0_combout ) # ((\prif.dataScr_wb [0] & (\prif.dataScr_wb [1] & \prif.pc_wb [11])))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.pc_wb [11]),
	.datad(\Mux153~0_combout ),
	.cin(gnd),
	.combout(\Mux153~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux153~1 .lut_mask = 16'hFF80;
defparam \Mux153~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N16
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (!ptBScr & ((always01 & ((\Mux153~1_combout ))) # (!always01 & (\prif.rdat2_ex [11]))))

	.dataa(\prif.rdat2_ex [11]),
	.datab(\Mux153~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'h00CA;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N30
cycloneive_lcell_comb \Mux84~2 (
// Equation(s):
// \Mux84~2_combout  = (\Mux52~0_combout ) # ((prifdmemaddr_11 & (ptBScr & !always01)))

	.dataa(prifdmemaddr_11),
	.datab(\HU|ptBScr~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux52~0_combout ),
	.cin(gnd),
	.combout(\Mux84~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux84~2 .lut_mask = 16'hFF08;
defparam \Mux84~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y26_N9
dffeas \prif.dmemload_wb[10] (
	.clk(CLK),
	.d(\PR|dmemload_wb~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[10] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y26_N31
dffeas \prif.dmemaddr_wb[10] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[10] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N16
cycloneive_lcell_comb \Mux154~0 (
// Equation(s):
// \Mux154~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [10]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [10]))))

	.dataa(\prif.dmemaddr_wb [10]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.dmemload_wb [10]),
	.datad(\prif.dataScr_wb [1]),
	.cin(gnd),
	.combout(\Mux154~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux154~0 .lut_mask = 16'h00E2;
defparam \Mux154~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y26_N23
dffeas \prif.pc_wb[10] (
	.clk(CLK),
	.d(\PR|pc_wb~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[10] .is_wysiwyg = "true";
defparam \prif.pc_wb[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N24
cycloneive_lcell_comb \Mux154~1 (
// Equation(s):
// \Mux154~1_combout  = (\Mux154~0_combout ) # ((\prif.pc_wb [10] & (\prif.dataScr_wb [0] & \prif.dataScr_wb [1])))

	.dataa(\prif.pc_wb [10]),
	.datab(\Mux154~0_combout ),
	.datac(\prif.dataScr_wb [0]),
	.datad(\prif.dataScr_wb [1]),
	.cin(gnd),
	.combout(\Mux154~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux154~1 .lut_mask = 16'hECCC;
defparam \Mux154~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N18
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (!ptBScr & ((always01 & (\Mux154~1_combout )) # (!always01 & ((\prif.rdat2_ex [10])))))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(\Mux154~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\prif.rdat2_ex [10]),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'h4540;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N12
cycloneive_lcell_comb \Mux85~2 (
// Equation(s):
// \Mux85~2_combout  = (\Mux53~0_combout ) # ((ptBScr & (prifdmemaddr_10 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_10),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux53~0_combout ),
	.cin(gnd),
	.combout(\Mux85~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux85~2 .lut_mask = 16'hFF08;
defparam \Mux85~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y28_N29
dffeas \prif.dmemload_wb[9] (
	.clk(CLK),
	.d(\PR|dmemload_wb~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[9] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y28_N7
dffeas \prif.dmemaddr_wb[9] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[9] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N16
cycloneive_lcell_comb \Mux155~0 (
// Equation(s):
// \Mux155~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [9]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [9]))))

	.dataa(\prif.dmemaddr_wb [9]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dmemload_wb [9]),
	.cin(gnd),
	.combout(\Mux155~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux155~0 .lut_mask = 16'h0E02;
defparam \Mux155~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N23
dffeas \prif.pc_wb[9] (
	.clk(CLK),
	.d(\PR|pc_wb~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[9] .is_wysiwyg = "true";
defparam \prif.pc_wb[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N22
cycloneive_lcell_comb \Mux155~1 (
// Equation(s):
// \Mux155~1_combout  = (\Mux155~0_combout ) # ((\prif.dataScr_wb [1] & (\prif.pc_wb [9] & \prif.dataScr_wb [0])))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.pc_wb [9]),
	.datac(\prif.dataScr_wb [0]),
	.datad(\Mux155~0_combout ),
	.cin(gnd),
	.combout(\Mux155~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux155~1 .lut_mask = 16'hFF80;
defparam \Mux155~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N20
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (!ptBScr & ((always01 & ((\Mux155~1_combout ))) # (!always01 & (\prif.rdat2_ex [9]))))

	.dataa(\HU|always0~5_combout ),
	.datab(\prif.rdat2_ex [9]),
	.datac(\Mux155~1_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'h00E4;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N30
cycloneive_lcell_comb \Mux86~2 (
// Equation(s):
// \Mux86~2_combout  = (\Mux54~0_combout ) # ((!always01 & (prifdmemaddr_9 & ptBScr)))

	.dataa(\HU|always0~5_combout ),
	.datab(prifdmemaddr_9),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\Mux54~0_combout ),
	.cin(gnd),
	.combout(\Mux86~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux86~2 .lut_mask = 16'hFF40;
defparam \Mux86~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y28_N3
dffeas \prif.dmemload_wb[6] (
	.clk(CLK),
	.d(\PR|dmemload_wb~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[6] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N15
dffeas \prif.dmemaddr_wb[6] (
	.clk(CLK),
	.d(gnd),
	.asdata(\PR|dmemaddr_wb~16_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[6] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N14
cycloneive_lcell_comb \Mux158~0 (
// Equation(s):
// \Mux158~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [6])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [6])))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dmemload_wb [6]),
	.datac(\prif.dmemaddr_wb [6]),
	.datad(\prif.dataScr_wb [1]),
	.cin(gnd),
	.combout(\Mux158~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux158~0 .lut_mask = 16'h00D8;
defparam \Mux158~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N25
dffeas \prif.pc_wb[6] (
	.clk(CLK),
	.d(\PR|pc_wb~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[6] .is_wysiwyg = "true";
defparam \prif.pc_wb[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N20
cycloneive_lcell_comb \Mux158~1 (
// Equation(s):
// \Mux158~1_combout  = (\Mux158~0_combout ) # ((\prif.dataScr_wb [0] & (\prif.dataScr_wb [1] & \prif.pc_wb [6])))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\Mux158~0_combout ),
	.datad(\prif.pc_wb [6]),
	.cin(gnd),
	.combout(\Mux158~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux158~1 .lut_mask = 16'hF8F0;
defparam \Mux158~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N2
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (!ptBScr & ((always01 & ((\Mux158~1_combout ))) # (!always01 & (\prif.rdat2_ex [6]))))

	.dataa(\prif.rdat2_ex [6]),
	.datab(\Mux158~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'h00CA;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N20
cycloneive_lcell_comb \Mux89~3 (
// Equation(s):
// \Mux89~3_combout  = (\Mux57~0_combout ) # ((ptBScr & (prifdmemaddr_6 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_6),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux57~0_combout ),
	.cin(gnd),
	.combout(\Mux89~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux89~3 .lut_mask = 16'hFF08;
defparam \Mux89~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y26_N17
dffeas \prif.dmemload_wb[27] (
	.clk(CLK),
	.d(\PR|dmemload_wb~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[27] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y26_N11
dffeas \prif.imm_wb[11] (
	.clk(CLK),
	.d(\PR|imm_wb~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[11] .is_wysiwyg = "true";
defparam \prif.imm_wb[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y26_N1
dffeas \prif.dmemaddr_wb[27] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[27] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N18
cycloneive_lcell_comb \Mux137~0 (
// Equation(s):
// \Mux137~0_combout  = (\prif.dataScr_wb [1] & ((\prif.imm_wb [11]) # ((\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & (((!\prif.dataScr_wb [0] & \prif.dmemaddr_wb [27]))))

	.dataa(\prif.imm_wb [11]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dataScr_wb [0]),
	.datad(\prif.dmemaddr_wb [27]),
	.cin(gnd),
	.combout(\Mux137~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux137~0 .lut_mask = 16'hCBC8;
defparam \Mux137~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y26_N13
dffeas \prif.pc_wb[27] (
	.clk(CLK),
	.d(\PR|pc_wb~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[27] .is_wysiwyg = "true";
defparam \prif.pc_wb[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N22
cycloneive_lcell_comb \Mux137~1 (
// Equation(s):
// \Mux137~1_combout  = (\prif.dataScr_wb [0] & ((\Mux137~0_combout  & (\prif.pc_wb [27])) # (!\Mux137~0_combout  & ((\prif.dmemload_wb [27]))))) # (!\prif.dataScr_wb [0] & (((\Mux137~0_combout ))))

	.dataa(\prif.pc_wb [27]),
	.datab(\prif.dmemload_wb [27]),
	.datac(\prif.dataScr_wb [0]),
	.datad(\Mux137~0_combout ),
	.cin(gnd),
	.combout(\Mux137~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux137~1 .lut_mask = 16'hAFC0;
defparam \Mux137~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N24
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (ptBScr & (((always01) # (prifdmemaddr_27)))) # (!ptBScr & (\prif.rdat2_ex [27] & (!always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(\prif.rdat2_ex [27]),
	.datac(\HU|always0~5_combout ),
	.datad(prifdmemaddr_27),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hAEA4;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N6
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (always01 & ((\Mux36~0_combout  & (\prif.imm_mem [11])) # (!\Mux36~0_combout  & ((\Mux137~1_combout ))))) # (!always01 & (((\Mux36~0_combout ))))

	.dataa(\prif.imm_mem [11]),
	.datab(\HU|always0~5_combout ),
	.datac(\Mux137~1_combout ),
	.datad(\Mux36~0_combout ),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hBBC0;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N20
cycloneive_lcell_comb \Mux68~0 (
// Equation(s):
// \Mux68~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux36~1_combout )))))

	.dataa(\prif.instr_ex [15]),
	.datab(\prif.ALUScr_ex [1]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux36~1_combout ),
	.cin(gnd),
	.combout(\Mux68~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux68~0 .lut_mask = 16'h2320;
defparam \Mux68~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y27_N5
dffeas \prif.dmemload_wb[23] (
	.clk(CLK),
	.d(\PR|dmemload_wb~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[23] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y27_N15
dffeas \prif.imm_wb[7] (
	.clk(CLK),
	.d(\PR|imm_wb~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[7] .is_wysiwyg = "true";
defparam \prif.imm_wb[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y27_N25
dffeas \prif.dmemaddr_wb[23] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[23] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N18
cycloneive_lcell_comb \Mux141~0 (
// Equation(s):
// \Mux141~0_combout  = (\prif.dataScr_wb [1] & (((\prif.imm_wb [7]) # (\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & (\prif.dmemaddr_wb [23] & ((!\prif.dataScr_wb [0]))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dmemaddr_wb [23]),
	.datac(\prif.imm_wb [7]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux141~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux141~0 .lut_mask = 16'hAAE4;
defparam \Mux141~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y27_N13
dffeas \prif.pc_wb[23] (
	.clk(CLK),
	.d(\PR|pc_wb~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[23] .is_wysiwyg = "true";
defparam \prif.pc_wb[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N10
cycloneive_lcell_comb \Mux141~1 (
// Equation(s):
// \Mux141~1_combout  = (\Mux141~0_combout  & ((\prif.pc_wb [23]) # ((!\prif.dataScr_wb [0])))) # (!\Mux141~0_combout  & (((\prif.dmemload_wb [23] & \prif.dataScr_wb [0]))))

	.dataa(\prif.pc_wb [23]),
	.datab(\Mux141~0_combout ),
	.datac(\prif.dmemload_wb [23]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux141~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux141~1 .lut_mask = 16'hB8CC;
defparam \Mux141~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N10
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (ptBScr & (((prifdmemaddr_23) # (always01)))) # (!ptBScr & (\prif.rdat2_ex [23] & ((!always01))))

	.dataa(\prif.rdat2_ex [23]),
	.datab(\HU|ptBScr~1_combout ),
	.datac(prifdmemaddr_23),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hCCE2;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N24
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (\Mux40~0_combout  & ((\prif.imm_mem [7]) # ((!always01)))) # (!\Mux40~0_combout  & (((\Mux141~1_combout  & always01))))

	.dataa(\Mux40~0_combout ),
	.datab(\prif.imm_mem [7]),
	.datac(\Mux141~1_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hD8AA;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N26
cycloneive_lcell_comb \Mux72~0 (
// Equation(s):
// \Mux72~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux40~1_combout )))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.instr_ex [15]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux40~1_combout ),
	.cin(gnd),
	.combout(\Mux72~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux72~0 .lut_mask = 16'h4540;
defparam \Mux72~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y29_N19
dffeas \prif.imm_wb[2] (
	.clk(CLK),
	.d(\PR|imm_wb~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[2] .is_wysiwyg = "true";
defparam \prif.imm_wb[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N1
dffeas \prif.dmemload_wb[18] (
	.clk(CLK),
	.d(\PR|dmemload_wb~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[18] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y29_N3
dffeas \prif.dmemaddr_wb[18] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[18] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N28
cycloneive_lcell_comb \Mux146~0 (
// Equation(s):
// \Mux146~0_combout  = (\prif.dataScr_wb [0] & ((\prif.dmemload_wb [18]) # ((\prif.dataScr_wb [1])))) # (!\prif.dataScr_wb [0] & (((!\prif.dataScr_wb [1] & \prif.dmemaddr_wb [18]))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dmemload_wb [18]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dmemaddr_wb [18]),
	.cin(gnd),
	.combout(\Mux146~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux146~0 .lut_mask = 16'hADA8;
defparam \Mux146~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y29_N31
dffeas \prif.pc_wb[18] (
	.clk(CLK),
	.d(\PR|pc_wb~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[18] .is_wysiwyg = "true";
defparam \prif.pc_wb[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N24
cycloneive_lcell_comb \Mux146~1 (
// Equation(s):
// \Mux146~1_combout  = (\prif.dataScr_wb [1] & ((\Mux146~0_combout  & ((\prif.pc_wb [18]))) # (!\Mux146~0_combout  & (\prif.imm_wb [2])))) # (!\prif.dataScr_wb [1] & (((\Mux146~0_combout ))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.imm_wb [2]),
	.datac(\prif.pc_wb [18]),
	.datad(\Mux146~0_combout ),
	.cin(gnd),
	.combout(\Mux146~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux146~1 .lut_mask = 16'hF588;
defparam \Mux146~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N10
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (always01 & (((ptBScr) # (\Mux146~1_combout )))) # (!always01 & (\prif.rdat2_ex [18] & (!ptBScr)))

	.dataa(\HU|always0~5_combout ),
	.datab(\prif.rdat2_ex [18]),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\Mux146~1_combout ),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hAEA4;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N12
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (ptBScr & ((\Mux45~0_combout  & ((\prif.imm_mem [2]))) # (!\Mux45~0_combout  & (prifdmemaddr_18)))) # (!ptBScr & (((\Mux45~0_combout ))))

	.dataa(prifdmemaddr_18),
	.datab(\prif.imm_mem [2]),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\Mux45~0_combout ),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hCFA0;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N14
cycloneive_lcell_comb \Mux77~0 (
// Equation(s):
// \Mux77~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux45~1_combout )))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.instr_ex [15]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux45~1_combout ),
	.cin(gnd),
	.combout(\Mux77~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux77~0 .lut_mask = 16'h4540;
defparam \Mux77~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y27_N27
dffeas \prif.imm_wb[8] (
	.clk(CLK),
	.d(\PR|imm_wb~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[8] .is_wysiwyg = "true";
defparam \prif.imm_wb[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N17
dffeas \prif.dmemload_wb[24] (
	.clk(CLK),
	.d(\PR|dmemload_wb~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[24] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N23
dffeas \prif.dmemaddr_wb[24] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[24] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N20
cycloneive_lcell_comb \Mux140~0 (
// Equation(s):
// \Mux140~0_combout  = (\prif.dataScr_wb [1] & (((\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [24]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [24]))))

	.dataa(\prif.dmemaddr_wb [24]),
	.datab(\prif.dmemload_wb [24]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux140~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux140~0 .lut_mask = 16'hFC0A;
defparam \Mux140~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y27_N19
dffeas \prif.pc_wb[24] (
	.clk(CLK),
	.d(\PR|pc_wb~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[24] .is_wysiwyg = "true";
defparam \prif.pc_wb[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N28
cycloneive_lcell_comb \Mux140~1 (
// Equation(s):
// \Mux140~1_combout  = (\prif.dataScr_wb [1] & ((\Mux140~0_combout  & (\prif.pc_wb [24])) # (!\Mux140~0_combout  & ((\prif.imm_wb [8]))))) # (!\prif.dataScr_wb [1] & (((\Mux140~0_combout ))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.pc_wb [24]),
	.datac(\prif.imm_wb [8]),
	.datad(\Mux140~0_combout ),
	.cin(gnd),
	.combout(\Mux140~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux140~1 .lut_mask = 16'hDDA0;
defparam \Mux140~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N14
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (ptBScr & (((always01)))) # (!ptBScr & ((always01 & ((\Mux140~1_combout ))) # (!always01 & (\prif.rdat2_ex [24]))))

	.dataa(\prif.rdat2_ex [24]),
	.datab(\Mux140~1_combout ),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hFC0A;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N24
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (ptBScr & ((\Mux39~0_combout  & (\prif.imm_mem [8])) # (!\Mux39~0_combout  & ((prifdmemaddr_24))))) # (!ptBScr & (((\Mux39~0_combout ))))

	.dataa(\prif.imm_mem [8]),
	.datab(\HU|ptBScr~1_combout ),
	.datac(\Mux39~0_combout ),
	.datad(prifdmemaddr_24),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hBCB0;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N30
cycloneive_lcell_comb \Mux71~0 (
// Equation(s):
// \Mux71~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux39~1_combout )))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.instr_ex [15]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux39~1_combout ),
	.cin(gnd),
	.combout(\Mux71~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux71~0 .lut_mask = 16'h4540;
defparam \Mux71~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y27_N1
dffeas \prif.imm_wb[0] (
	.clk(CLK),
	.d(\PR|imm_wb~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[0] .is_wysiwyg = "true";
defparam \prif.imm_wb[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N5
dffeas \prif.dmemload_wb[16] (
	.clk(CLK),
	.d(\PR|dmemload_wb~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[16] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N27
dffeas \prif.dmemaddr_wb[16] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[16] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N8
cycloneive_lcell_comb \Mux148~0 (
// Equation(s):
// \Mux148~0_combout  = (\prif.dataScr_wb [1] & (((\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [16])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [16])))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dmemload_wb [16]),
	.datac(\prif.dmemaddr_wb [16]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux148~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux148~0 .lut_mask = 16'hEE50;
defparam \Mux148~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y27_N3
dffeas \prif.pc_wb[16] (
	.clk(CLK),
	.d(\PR|pc_wb~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[16] .is_wysiwyg = "true";
defparam \prif.pc_wb[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N16
cycloneive_lcell_comb \Mux148~1 (
// Equation(s):
// \Mux148~1_combout  = (\prif.dataScr_wb [1] & ((\Mux148~0_combout  & ((\prif.pc_wb [16]))) # (!\Mux148~0_combout  & (\prif.imm_wb [0])))) # (!\prif.dataScr_wb [1] & (((\Mux148~0_combout ))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.imm_wb [0]),
	.datac(\Mux148~0_combout ),
	.datad(\prif.pc_wb [16]),
	.cin(gnd),
	.combout(\Mux148~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux148~1 .lut_mask = 16'hF858;
defparam \Mux148~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N26
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (ptBScr & (always01)) # (!ptBScr & ((always01 & ((\Mux148~1_combout ))) # (!always01 & (\prif.rdat2_ex [16]))))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(\prif.rdat2_ex [16]),
	.datad(\Mux148~1_combout ),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hDC98;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N28
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (\Mux47~0_combout  & ((\prif.imm_mem [0]) # ((!ptBScr)))) # (!\Mux47~0_combout  & (((prifdmemaddr_16 & ptBScr))))

	.dataa(\prif.imm_mem [0]),
	.datab(prifdmemaddr_16),
	.datac(\Mux47~0_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hACF0;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N6
cycloneive_lcell_comb \Mux79~0 (
// Equation(s):
// \Mux79~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux47~1_combout )))))

	.dataa(\prif.instr_ex [15]),
	.datab(\prif.ALUScr_ex [1]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux47~1_combout ),
	.cin(gnd),
	.combout(\Mux79~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux79~0 .lut_mask = 16'h2320;
defparam \Mux79~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N9
dffeas \prif.dmemload_wb[19] (
	.clk(CLK),
	.d(\PR|dmemload_wb~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[19] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N23
dffeas \prif.imm_wb[3] (
	.clk(CLK),
	.d(\PR|imm_wb~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[3] .is_wysiwyg = "true";
defparam \prif.imm_wb[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N21
dffeas \prif.dmemaddr_wb[19] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[19] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N2
cycloneive_lcell_comb \Mux145~0 (
// Equation(s):
// \Mux145~0_combout  = (\prif.dataScr_wb [1] & ((\prif.imm_wb [3]) # ((\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & (((\prif.dmemaddr_wb [19] & !\prif.dataScr_wb [0]))))

	.dataa(\prif.imm_wb [3]),
	.datab(\prif.dmemaddr_wb [19]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux145~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux145~0 .lut_mask = 16'hF0AC;
defparam \Mux145~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y29_N17
dffeas \prif.pc_wb[19] (
	.clk(CLK),
	.d(\PR|pc_wb~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[19] .is_wysiwyg = "true";
defparam \prif.pc_wb[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N18
cycloneive_lcell_comb \Mux145~1 (
// Equation(s):
// \Mux145~1_combout  = (\prif.dataScr_wb [0] & ((\Mux145~0_combout  & (\prif.pc_wb [19])) # (!\Mux145~0_combout  & ((\prif.dmemload_wb [19]))))) # (!\prif.dataScr_wb [0] & (((\Mux145~0_combout ))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.pc_wb [19]),
	.datac(\prif.dmemload_wb [19]),
	.datad(\Mux145~0_combout ),
	.cin(gnd),
	.combout(\Mux145~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux145~1 .lut_mask = 16'hDDA0;
defparam \Mux145~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N12
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (ptBScr & (((prifdmemaddr_19) # (always01)))) # (!ptBScr & (\prif.rdat2_ex [19] & ((!always01))))

	.dataa(\prif.rdat2_ex [19]),
	.datab(prifdmemaddr_19),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hF0CA;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N6
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (\Mux44~0_combout  & (((\prif.imm_mem [3]) # (!always01)))) # (!\Mux44~0_combout  & (\Mux145~1_combout  & ((always01))))

	.dataa(\Mux44~0_combout ),
	.datab(\Mux145~1_combout ),
	.datac(\prif.imm_mem [3]),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hE4AA;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N14
cycloneive_lcell_comb \Mux76~0 (
// Equation(s):
// \Mux76~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & ((\prif.instr_ex [15]))) # (!\prif.ALUScr_ex [0] & (\Mux44~1_combout ))))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.ALUScr_ex [1]),
	.datac(\Mux44~1_combout ),
	.datad(\prif.instr_ex [15]),
	.cin(gnd),
	.combout(\Mux76~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux76~0 .lut_mask = 16'h3210;
defparam \Mux76~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y29_N19
dffeas \prif.dmemload_wb[17] (
	.clk(CLK),
	.d(\PR|dmemload_wb~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[17] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N1
dffeas \prif.imm_wb[1] (
	.clk(CLK),
	.d(\PR|imm_wb~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[1] .is_wysiwyg = "true";
defparam \prif.imm_wb[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N23
dffeas \prif.dmemaddr_wb[17] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[17] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N20
cycloneive_lcell_comb \Mux147~0 (
// Equation(s):
// \Mux147~0_combout  = (\prif.dataScr_wb [1] & (((\prif.imm_wb [1]) # (\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & (\prif.dmemaddr_wb [17] & ((!\prif.dataScr_wb [0]))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dmemaddr_wb [17]),
	.datac(\prif.imm_wb [1]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux147~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux147~0 .lut_mask = 16'hAAE4;
defparam \Mux147~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y28_N23
dffeas \prif.pc_wb[17] (
	.clk(CLK),
	.d(\PR|pc_wb~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[17] .is_wysiwyg = "true";
defparam \prif.pc_wb[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N14
cycloneive_lcell_comb \Mux147~1 (
// Equation(s):
// \Mux147~1_combout  = (\Mux147~0_combout  & ((\prif.pc_wb [17]) # ((!\prif.dataScr_wb [0])))) # (!\Mux147~0_combout  & (((\prif.dataScr_wb [0] & \prif.dmemload_wb [17]))))

	.dataa(\prif.pc_wb [17]),
	.datab(\Mux147~0_combout ),
	.datac(\prif.dataScr_wb [0]),
	.datad(\prif.dmemload_wb [17]),
	.cin(gnd),
	.combout(\Mux147~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux147~1 .lut_mask = 16'hBC8C;
defparam \Mux147~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N4
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (always01 & (((ptBScr)))) # (!always01 & ((ptBScr & ((prifdmemaddr_17))) # (!ptBScr & (\prif.rdat2_ex [17]))))

	.dataa(\HU|always0~5_combout ),
	.datab(\prif.rdat2_ex [17]),
	.datac(prifdmemaddr_17),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hFA44;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N12
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (\Mux46~0_combout  & ((\prif.imm_mem [1]) # ((!always01)))) # (!\Mux46~0_combout  & (((\Mux147~1_combout  & always01))))

	.dataa(\prif.imm_mem [1]),
	.datab(\Mux147~1_combout ),
	.datac(\Mux46~0_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hACF0;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N10
cycloneive_lcell_comb \Mux78~0 (
// Equation(s):
// \Mux78~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux46~1_combout )))))

	.dataa(\prif.instr_ex [15]),
	.datab(\prif.ALUScr_ex [1]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux46~1_combout ),
	.cin(gnd),
	.combout(\Mux78~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux78~0 .lut_mask = 16'h2320;
defparam \Mux78~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N21
dffeas \prif.dmemload_wb[21] (
	.clk(CLK),
	.d(\PR|dmemload_wb~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[21] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N1
dffeas \prif.imm_wb[5] (
	.clk(CLK),
	.d(\PR|imm_wb~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[5] .is_wysiwyg = "true";
defparam \prif.imm_wb[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N27
dffeas \prif.dmemaddr_wb[21] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[21] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N12
cycloneive_lcell_comb \Mux143~0 (
// Equation(s):
// \Mux143~0_combout  = (\prif.dataScr_wb [1] & (((\prif.imm_wb [5]) # (\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & (\prif.dmemaddr_wb [21] & ((!\prif.dataScr_wb [0]))))

	.dataa(\prif.dmemaddr_wb [21]),
	.datab(\prif.imm_wb [5]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux143~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux143~0 .lut_mask = 16'hF0CA;
defparam \Mux143~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y29_N19
dffeas \prif.pc_wb[21] (
	.clk(CLK),
	.d(\PR|pc_wb~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[21] .is_wysiwyg = "true";
defparam \prif.pc_wb[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N24
cycloneive_lcell_comb \Mux143~1 (
// Equation(s):
// \Mux143~1_combout  = (\prif.dataScr_wb [0] & ((\Mux143~0_combout  & (\prif.pc_wb [21])) # (!\Mux143~0_combout  & ((\prif.dmemload_wb [21]))))) # (!\prif.dataScr_wb [0] & (((\Mux143~0_combout ))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.pc_wb [21]),
	.datac(\prif.dmemload_wb [21]),
	.datad(\Mux143~0_combout ),
	.cin(gnd),
	.combout(\Mux143~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux143~1 .lut_mask = 16'hDDA0;
defparam \Mux143~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N14
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (ptBScr & (((prifdmemaddr_21) # (always01)))) # (!ptBScr & (\prif.rdat2_ex [21] & ((!always01))))

	.dataa(\prif.rdat2_ex [21]),
	.datab(prifdmemaddr_21),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hF0CA;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N20
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (\Mux42~0_combout  & (((\prif.imm_mem [5])) # (!always01))) # (!\Mux42~0_combout  & (always01 & ((\Mux143~1_combout ))))

	.dataa(\Mux42~0_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(\prif.imm_mem [5]),
	.datad(\Mux143~1_combout ),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hE6A2;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N30
cycloneive_lcell_comb \Mux74~0 (
// Equation(s):
// \Mux74~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux42~1_combout )))))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.instr_ex [15]),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\Mux42~1_combout ),
	.cin(gnd),
	.combout(\Mux74~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux74~0 .lut_mask = 16'h0D08;
defparam \Mux74~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N27
dffeas \prif.imm_wb[4] (
	.clk(CLK),
	.d(\PR|imm_wb~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[4] .is_wysiwyg = "true";
defparam \prif.imm_wb[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N13
dffeas \prif.dmemload_wb[20] (
	.clk(CLK),
	.d(\PR|dmemload_wb~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[20] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N19
dffeas \prif.dmemaddr_wb[20] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[20] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N28
cycloneive_lcell_comb \Mux144~0 (
// Equation(s):
// \Mux144~0_combout  = (\prif.dataScr_wb [0] & ((\prif.dmemload_wb [20]) # ((\prif.dataScr_wb [1])))) # (!\prif.dataScr_wb [0] & (((!\prif.dataScr_wb [1] & \prif.dmemaddr_wb [20]))))

	.dataa(\prif.dmemload_wb [20]),
	.datab(\prif.dataScr_wb [0]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dmemaddr_wb [20]),
	.cin(gnd),
	.combout(\Mux144~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux144~0 .lut_mask = 16'hCBC8;
defparam \Mux144~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y31_N31
dffeas \prif.pc_wb[20] (
	.clk(CLK),
	.d(\PR|pc_wb~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[20] .is_wysiwyg = "true";
defparam \prif.pc_wb[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N8
cycloneive_lcell_comb \Mux144~1 (
// Equation(s):
// \Mux144~1_combout  = (\prif.dataScr_wb [1] & ((\Mux144~0_combout  & ((\prif.pc_wb [20]))) # (!\Mux144~0_combout  & (\prif.imm_wb [4])))) # (!\prif.dataScr_wb [1] & (((\Mux144~0_combout ))))

	.dataa(\prif.imm_wb [4]),
	.datab(\prif.pc_wb [20]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\Mux144~0_combout ),
	.cin(gnd),
	.combout(\Mux144~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux144~1 .lut_mask = 16'hCFA0;
defparam \Mux144~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N2
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (ptBScr & (((always01)))) # (!ptBScr & ((always01 & (\Mux144~1_combout )) # (!always01 & ((\prif.rdat2_ex [20])))))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(\Mux144~1_combout ),
	.datac(\prif.rdat2_ex [20]),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hEE50;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N20
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (\Mux43~0_combout  & ((\prif.imm_mem [4]) # ((!ptBScr)))) # (!\Mux43~0_combout  & (((prifdmemaddr_20 & ptBScr))))

	.dataa(\prif.imm_mem [4]),
	.datab(\Mux43~0_combout ),
	.datac(prifdmemaddr_20),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hB8CC;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N20
cycloneive_lcell_comb \Mux75~0 (
// Equation(s):
// \Mux75~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux43~1_combout )))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.ALUScr_ex [0]),
	.datac(\prif.instr_ex [15]),
	.datad(\Mux43~1_combout ),
	.cin(gnd),
	.combout(\Mux75~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux75~0 .lut_mask = 16'h5140;
defparam \Mux75~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y26_N1
dffeas \prif.imm_wb[12] (
	.clk(CLK),
	.d(\PR|imm_wb~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[12] .is_wysiwyg = "true";
defparam \prif.imm_wb[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y26_N23
dffeas \prif.dmemload_wb[28] (
	.clk(CLK),
	.d(\PR|dmemload_wb~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[28] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y26_N5
dffeas \prif.dmemaddr_wb[28] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[28] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N26
cycloneive_lcell_comb \Mux136~0 (
// Equation(s):
// \Mux136~0_combout  = (\prif.dataScr_wb [1] & (((\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [28])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [28])))))

	.dataa(\prif.dmemload_wb [28]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dmemaddr_wb [28]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux136~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux136~0 .lut_mask = 16'hEE30;
defparam \Mux136~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y26_N13
dffeas \prif.pc_wb[28] (
	.clk(CLK),
	.d(\PR|pc_wb~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[28] .is_wysiwyg = "true";
defparam \prif.pc_wb[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N2
cycloneive_lcell_comb \Mux136~1 (
// Equation(s):
// \Mux136~1_combout  = (\Mux136~0_combout  & ((\prif.pc_wb [28]) # ((!\prif.dataScr_wb [1])))) # (!\Mux136~0_combout  & (((\prif.imm_wb [12] & \prif.dataScr_wb [1]))))

	.dataa(\prif.pc_wb [28]),
	.datab(\prif.imm_wb [12]),
	.datac(\Mux136~0_combout ),
	.datad(\prif.dataScr_wb [1]),
	.cin(gnd),
	.combout(\Mux136~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux136~1 .lut_mask = 16'hACF0;
defparam \Mux136~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N28
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (always01 & (((ptBScr) # (\Mux136~1_combout )))) # (!always01 & (\prif.rdat2_ex [28] & (!ptBScr)))

	.dataa(\prif.rdat2_ex [28]),
	.datab(\HU|always0~5_combout ),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\Mux136~1_combout ),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hCEC2;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N10
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (ptBScr & ((\Mux35~0_combout  & (\prif.imm_mem [12])) # (!\Mux35~0_combout  & ((prifdmemaddr_28))))) # (!ptBScr & (((\Mux35~0_combout ))))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(\prif.imm_mem [12]),
	.datac(prifdmemaddr_28),
	.datad(\Mux35~0_combout ),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hDDA0;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N16
cycloneive_lcell_comb \Mux67~0 (
// Equation(s):
// \Mux67~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux35~1_combout )))))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.instr_ex [15]),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\Mux35~1_combout ),
	.cin(gnd),
	.combout(\Mux67~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux67~0 .lut_mask = 16'h0D08;
defparam \Mux67~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y27_N15
dffeas \prif.imm_wb[10] (
	.clk(CLK),
	.d(\PR|imm_wb~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[10] .is_wysiwyg = "true";
defparam \prif.imm_wb[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N29
dffeas \prif.dmemload_wb[26] (
	.clk(CLK),
	.d(\PR|dmemload_wb~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[26] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N11
dffeas \prif.dmemaddr_wb[26] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[26] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N8
cycloneive_lcell_comb \Mux138~0 (
// Equation(s):
// \Mux138~0_combout  = (\prif.dataScr_wb [1] & (((\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [26]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [26]))))

	.dataa(\prif.dmemaddr_wb [26]),
	.datab(\prif.dmemload_wb [26]),
	.datac(\prif.dataScr_wb [1]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux138~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux138~0 .lut_mask = 16'hFC0A;
defparam \Mux138~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y27_N7
dffeas \prif.pc_wb[26] (
	.clk(CLK),
	.d(\PR|pc_wb~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[26] .is_wysiwyg = "true";
defparam \prif.pc_wb[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N0
cycloneive_lcell_comb \Mux138~1 (
// Equation(s):
// \Mux138~1_combout  = (\prif.dataScr_wb [1] & ((\Mux138~0_combout  & ((\prif.pc_wb [26]))) # (!\Mux138~0_combout  & (\prif.imm_wb [10])))) # (!\prif.dataScr_wb [1] & (((\Mux138~0_combout ))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.imm_wb [10]),
	.datac(\Mux138~0_combout ),
	.datad(\prif.pc_wb [26]),
	.cin(gnd),
	.combout(\Mux138~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux138~1 .lut_mask = 16'hF858;
defparam \Mux138~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N22
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (ptBScr & (((always01)))) # (!ptBScr & ((always01 & ((\Mux138~1_combout ))) # (!always01 & (\prif.rdat2_ex [26]))))

	.dataa(\prif.rdat2_ex [26]),
	.datab(\HU|ptBScr~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux138~1_combout ),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hF2C2;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N24
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (\Mux37~0_combout  & ((\prif.imm_mem [10]) # ((!ptBScr)))) # (!\Mux37~0_combout  & (((ptBScr & prifdmemaddr_26))))

	.dataa(\Mux37~0_combout ),
	.datab(\prif.imm_mem [10]),
	.datac(\HU|ptBScr~1_combout ),
	.datad(prifdmemaddr_26),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hDA8A;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N30
cycloneive_lcell_comb \Mux69~0 (
// Equation(s):
// \Mux69~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux37~1_combout )))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.ALUScr_ex [0]),
	.datac(\prif.instr_ex [15]),
	.datad(\Mux37~1_combout ),
	.cin(gnd),
	.combout(\Mux69~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux69~0 .lut_mask = 16'h5140;
defparam \Mux69~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y30_N31
dffeas \prif.dmemload_wb[8] (
	.clk(CLK),
	.d(\PR|dmemload_wb~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[8] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N3
dffeas \prif.dmemaddr_wb[8] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[8] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N0
cycloneive_lcell_comb \Mux156~0 (
// Equation(s):
// \Mux156~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [8])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [8])))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dmemload_wb [8]),
	.datad(\prif.dmemaddr_wb [8]),
	.cin(gnd),
	.combout(\Mux156~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux156~0 .lut_mask = 16'h3120;
defparam \Mux156~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y29_N17
dffeas \prif.pc_wb[8] (
	.clk(CLK),
	.d(\PR|pc_wb~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[8] .is_wysiwyg = "true";
defparam \prif.pc_wb[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N22
cycloneive_lcell_comb \Mux156~1 (
// Equation(s):
// \Mux156~1_combout  = (\Mux156~0_combout ) # ((\prif.dataScr_wb [0] & (\prif.dataScr_wb [1] & \prif.pc_wb [8])))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.pc_wb [8]),
	.datad(\Mux156~0_combout ),
	.cin(gnd),
	.combout(\Mux156~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux156~1 .lut_mask = 16'hFF80;
defparam \Mux156~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N30
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (!ptBScr & ((always01 & ((\Mux156~1_combout ))) # (!always01 & (\prif.rdat2_ex [8]))))

	.dataa(\prif.rdat2_ex [8]),
	.datab(\HU|ptBScr~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux156~1_combout ),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'h3202;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N12
cycloneive_lcell_comb \Mux87~2 (
// Equation(s):
// \Mux87~2_combout  = (\Mux55~0_combout ) # ((!always01 & (ptBScr & prifdmemaddr_8)))

	.dataa(\Mux55~0_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(\HU|ptBScr~1_combout ),
	.datad(prifdmemaddr_8),
	.cin(gnd),
	.combout(\Mux87~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux87~2 .lut_mask = 16'hBAAA;
defparam \Mux87~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y29_N9
dffeas \prif.dmemload_wb[7] (
	.clk(CLK),
	.d(\PR|dmemload_wb~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[7] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N11
dffeas \prif.dmemaddr_wb[7] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[7] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N4
cycloneive_lcell_comb \Mux157~0 (
// Equation(s):
// \Mux157~0_combout  = (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & (\prif.dmemload_wb [7])) # (!\prif.dataScr_wb [0] & ((\prif.dmemaddr_wb [7])))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\prif.dmemload_wb [7]),
	.datad(\prif.dmemaddr_wb [7]),
	.cin(gnd),
	.combout(\Mux157~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux157~0 .lut_mask = 16'h3120;
defparam \Mux157~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y33_N19
dffeas \prif.pc_wb[7] (
	.clk(CLK),
	.d(\PR|pc_wb~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[7] .is_wysiwyg = "true";
defparam \prif.pc_wb[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N18
cycloneive_lcell_comb \Mux157~1 (
// Equation(s):
// \Mux157~1_combout  = (\Mux157~0_combout ) # ((\prif.dataScr_wb [0] & (\prif.dataScr_wb [1] & \prif.pc_wb [7])))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dataScr_wb [1]),
	.datac(\Mux157~0_combout ),
	.datad(\prif.pc_wb [7]),
	.cin(gnd),
	.combout(\Mux157~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux157~1 .lut_mask = 16'hF8F0;
defparam \Mux157~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N2
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (!ptBScr & ((always01 & (\Mux157~1_combout )) # (!always01 & ((\prif.rdat2_ex [7])))))

	.dataa(\Mux157~1_combout ),
	.datab(\HU|ptBScr~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\prif.rdat2_ex [7]),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'h2320;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N8
cycloneive_lcell_comb \Mux88~2 (
// Equation(s):
// \Mux88~2_combout  = (\Mux56~0_combout ) # ((ptBScr & (prifdmemaddr_7 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_7),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux56~0_combout ),
	.cin(gnd),
	.combout(\Mux88~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux88~2 .lut_mask = 16'hFF08;
defparam \Mux88~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y27_N9
dffeas \prif.imm_wb[6] (
	.clk(CLK),
	.d(\PR|imm_wb~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[6] .is_wysiwyg = "true";
defparam \prif.imm_wb[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y27_N31
dffeas \prif.dmemload_wb[22] (
	.clk(CLK),
	.d(\PR|dmemload_wb~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[22] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y27_N29
dffeas \prif.dmemaddr_wb[22] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[22] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N2
cycloneive_lcell_comb \Mux142~0 (
// Equation(s):
// \Mux142~0_combout  = (\prif.dataScr_wb [1] & (((\prif.dataScr_wb [0])))) # (!\prif.dataScr_wb [1] & ((\prif.dataScr_wb [0] & ((\prif.dmemload_wb [22]))) # (!\prif.dataScr_wb [0] & (\prif.dmemaddr_wb [22]))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.dmemaddr_wb [22]),
	.datac(\prif.dmemload_wb [22]),
	.datad(\prif.dataScr_wb [0]),
	.cin(gnd),
	.combout(\Mux142~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux142~0 .lut_mask = 16'hFA44;
defparam \Mux142~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y27_N21
dffeas \prif.pc_wb[22] (
	.clk(CLK),
	.d(\PR|pc_wb~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[22] .is_wysiwyg = "true";
defparam \prif.pc_wb[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N22
cycloneive_lcell_comb \Mux142~1 (
// Equation(s):
// \Mux142~1_combout  = (\prif.dataScr_wb [1] & ((\Mux142~0_combout  & (\prif.pc_wb [22])) # (!\Mux142~0_combout  & ((\prif.imm_wb [6]))))) # (!\prif.dataScr_wb [1] & (((\Mux142~0_combout ))))

	.dataa(\prif.dataScr_wb [1]),
	.datab(\prif.pc_wb [22]),
	.datac(\prif.imm_wb [6]),
	.datad(\Mux142~0_combout ),
	.cin(gnd),
	.combout(\Mux142~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux142~1 .lut_mask = 16'hDDA0;
defparam \Mux142~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N0
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (always01 & (((\Mux142~1_combout ) # (ptBScr)))) # (!always01 & (\prif.rdat2_ex [22] & ((!ptBScr))))

	.dataa(\prif.rdat2_ex [22]),
	.datab(\HU|always0~5_combout ),
	.datac(\Mux142~1_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hCCE2;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N2
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (ptBScr & ((\Mux41~0_combout  & (\prif.imm_mem [6])) # (!\Mux41~0_combout  & ((prifdmemaddr_22))))) # (!ptBScr & (((\Mux41~0_combout ))))

	.dataa(\prif.imm_mem [6]),
	.datab(\HU|ptBScr~1_combout ),
	.datac(prifdmemaddr_22),
	.datad(\Mux41~0_combout ),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hBBC0;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N8
cycloneive_lcell_comb \Mux73~0 (
// Equation(s):
// \Mux73~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux41~1_combout )))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.instr_ex [15]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux41~1_combout ),
	.cin(gnd),
	.combout(\Mux73~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux73~0 .lut_mask = 16'h4540;
defparam \Mux73~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y28_N13
dffeas \prif.dmemload_wb[25] (
	.clk(CLK),
	.d(\PR|dmemload_wb~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemload_wb [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemload_wb[25] .is_wysiwyg = "true";
defparam \prif.dmemload_wb[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N27
dffeas \prif.imm_wb[9] (
	.clk(CLK),
	.d(\PR|imm_wb~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.imm_wb [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.imm_wb[9] .is_wysiwyg = "true";
defparam \prif.imm_wb[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y28_N17
dffeas \prif.dmemaddr_wb[25] (
	.clk(CLK),
	.d(\PR|dmemaddr_wb~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.dmemaddr_wb [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr_wb[25] .is_wysiwyg = "true";
defparam \prif.dmemaddr_wb[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N14
cycloneive_lcell_comb \Mux139~0 (
// Equation(s):
// \Mux139~0_combout  = (\prif.dataScr_wb [0] & (((\prif.dataScr_wb [1])))) # (!\prif.dataScr_wb [0] & ((\prif.dataScr_wb [1] & ((\prif.imm_wb [9]))) # (!\prif.dataScr_wb [1] & (\prif.dmemaddr_wb [25]))))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\prif.dmemaddr_wb [25]),
	.datac(\prif.imm_wb [9]),
	.datad(\prif.dataScr_wb [1]),
	.cin(gnd),
	.combout(\Mux139~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux139~0 .lut_mask = 16'hFA44;
defparam \Mux139~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y28_N9
dffeas \prif.pc_wb[25] (
	.clk(CLK),
	.d(\PR|pc_wb~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_wb [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_wb[25] .is_wysiwyg = "true";
defparam \prif.pc_wb[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N6
cycloneive_lcell_comb \Mux139~1 (
// Equation(s):
// \Mux139~1_combout  = (\prif.dataScr_wb [0] & ((\Mux139~0_combout  & (\prif.pc_wb [25])) # (!\Mux139~0_combout  & ((\prif.dmemload_wb [25]))))) # (!\prif.dataScr_wb [0] & (\Mux139~0_combout ))

	.dataa(\prif.dataScr_wb [0]),
	.datab(\Mux139~0_combout ),
	.datac(\prif.pc_wb [25]),
	.datad(\prif.dmemload_wb [25]),
	.cin(gnd),
	.combout(\Mux139~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux139~1 .lut_mask = 16'hE6C4;
defparam \Mux139~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N4
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (always01 & (ptBScr)) # (!always01 & ((ptBScr & (prifdmemaddr_25)) # (!ptBScr & ((\prif.rdat2_ex [25])))))

	.dataa(\HU|always0~5_combout ),
	.datab(\HU|ptBScr~1_combout ),
	.datac(prifdmemaddr_25),
	.datad(\prif.rdat2_ex [25]),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hD9C8;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N2
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (\Mux38~0_combout  & (((\prif.imm_mem [9]) # (!always01)))) # (!\Mux38~0_combout  & (\Mux139~1_combout  & ((always01))))

	.dataa(\Mux139~1_combout ),
	.datab(\prif.imm_mem [9]),
	.datac(\Mux38~0_combout ),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hCAF0;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N0
cycloneive_lcell_comb \Mux70~0 (
// Equation(s):
// \Mux70~0_combout  = (!\prif.ALUScr_ex [1] & ((\prif.ALUScr_ex [0] & (\prif.instr_ex [15])) # (!\prif.ALUScr_ex [0] & ((\Mux38~1_combout )))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.instr_ex [15]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux38~1_combout ),
	.cin(gnd),
	.combout(\Mux70~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux70~0 .lut_mask = 16'h4540;
defparam \Mux70~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y30_N19
dffeas \prif.ALUOP_ex[2] (
	.clk(CLK),
	.d(\PR|ALUOP_ex~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.ALUOP_ex [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.ALUOP_ex[2] .is_wysiwyg = "true";
defparam \prif.ALUOP_ex[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y25_N31
dffeas \prif.ALUOP_ex[1] (
	.clk(CLK),
	.d(\PR|ALUOP_ex~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.ALUOP_ex [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.ALUOP_ex[1] .is_wysiwyg = "true";
defparam \prif.ALUOP_ex[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N24
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (always02 & (prifdmemaddr_2)) # (!always02 & ((\prif.rdat1_ex [2])))

	.dataa(prifdmemaddr_2),
	.datab(gnd),
	.datac(\prif.rdat1_ex [2]),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hAAF0;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N26
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (ptAScr & (\Mux162~1_combout  & ((!always02)))) # (!ptAScr & (((\Mux29~0_combout ))))

	.dataa(\Mux162~1_combout ),
	.datab(\Mux29~0_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'h0ACC;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N0
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (always02 & (prifdmemaddr_4)) # (!always02 & ((\prif.rdat1_ex [4])))

	.dataa(\HU|always0~6_combout ),
	.datab(gnd),
	.datac(prifdmemaddr_4),
	.datad(\prif.rdat1_ex [4]),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hF5A0;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N14
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (ptAScr & (\Mux160~1_combout  & ((!always02)))) # (!ptAScr & (((\Mux27~0_combout ))))

	.dataa(\Mux160~1_combout ),
	.datab(\Mux27~0_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'h0ACC;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N28
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (always02 & (prifdmemaddr_3)) # (!always02 & ((\prif.rdat1_ex [3])))

	.dataa(\HU|always0~6_combout ),
	.datab(gnd),
	.datac(prifdmemaddr_3),
	.datad(\prif.rdat1_ex [3]),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hF5A0;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N6
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (ptAScr & (((!always02 & \Mux161~1_combout )))) # (!ptAScr & (\Mux28~0_combout ))

	.dataa(\HU|ptAScr~4_combout ),
	.datab(\Mux28~0_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\Mux161~1_combout ),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'h4E44;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N2
cycloneive_lcell_comb \Mux93~1 (
// Equation(s):
// \Mux93~1_combout  = (ptBScr & (prifdmemaddr_2 & !always01))

	.dataa(gnd),
	.datab(\HU|ptBScr~1_combout ),
	.datac(prifdmemaddr_2),
	.datad(\HU|always0~5_combout ),
	.cin(gnd),
	.combout(\Mux93~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux93~1 .lut_mask = 16'h00C0;
defparam \Mux93~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N4
cycloneive_lcell_comb \Mux93~2 (
// Equation(s):
// \Mux93~2_combout  = (\Mux93~0_combout ) # ((\Mux89~2_combout  & ((\Mux61~0_combout ) # (\Mux93~1_combout ))))

	.dataa(\Mux93~0_combout ),
	.datab(\Mux61~0_combout ),
	.datac(\Mux89~2_combout ),
	.datad(\Mux93~1_combout ),
	.cin(gnd),
	.combout(\Mux93~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux93~2 .lut_mask = 16'hFAEA;
defparam \Mux93~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N18
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (always02 & ((prifdmemaddr_8))) # (!always02 & (\prif.rdat1_ex [8]))

	.dataa(gnd),
	.datab(\prif.rdat1_ex [8]),
	.datac(prifdmemaddr_8),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hF0CC;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N16
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (ptAScr & (\Mux156~1_combout  & ((!always02)))) # (!ptAScr & (((\Mux23~0_combout ))))

	.dataa(\Mux156~1_combout ),
	.datab(\Mux23~0_combout ),
	.datac(\HU|ptAScr~4_combout ),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'h0CAC;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N4
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (always02 & (prifdmemaddr_7)) # (!always02 & ((\prif.rdat1_ex [7])))

	.dataa(prifdmemaddr_7),
	.datab(gnd),
	.datac(\prif.rdat1_ex [7]),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hAAF0;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N6
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (ptAScr & (\Mux157~1_combout  & ((!always02)))) # (!ptAScr & (((\Mux24~0_combout ))))

	.dataa(\Mux157~1_combout ),
	.datab(\HU|ptAScr~4_combout ),
	.datac(\Mux24~0_combout ),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'h30B8;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N26
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (always02 & (prifdmemaddr_6)) # (!always02 & ((\prif.rdat1_ex [6])))

	.dataa(gnd),
	.datab(prifdmemaddr_6),
	.datac(\HU|always0~6_combout ),
	.datad(\prif.rdat1_ex [6]),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hCFC0;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N8
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (ptAScr & (((\Mux158~1_combout  & !always02)))) # (!ptAScr & (\Mux25~0_combout ))

	.dataa(\Mux25~0_combout ),
	.datab(\Mux158~1_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'h0CAA;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N0
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (always02 & ((prifdmemaddr_5))) # (!always02 & (\prif.rdat1_ex [5]))

	.dataa(gnd),
	.datab(\prif.rdat1_ex [5]),
	.datac(\HU|always0~6_combout ),
	.datad(prifdmemaddr_5),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hFC0C;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N30
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (ptAScr & (\Mux159~1_combout  & (!always02))) # (!ptAScr & (((\Mux26~0_combout ))))

	.dataa(\HU|ptAScr~4_combout ),
	.datab(\Mux159~1_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\Mux26~0_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'h5D08;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N24
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (always02 & ((ptAScr & (\prif.imm_mem [0])) # (!ptAScr & ((prifdmemaddr_16))))) # (!always02 & (((ptAScr))))

	.dataa(\prif.imm_mem [0]),
	.datab(prifdmemaddr_16),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hAFC0;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N30
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (always02 & (((\Mux15~0_combout )))) # (!always02 & ((\Mux15~0_combout  & ((\Mux148~1_combout ))) # (!\Mux15~0_combout  & (\prif.rdat1_ex [16]))))

	.dataa(\prif.rdat1_ex [16]),
	.datab(\Mux148~1_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hFC0A;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N4
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (always02 & ((prifdmemaddr_15))) # (!always02 & (\prif.rdat1_ex [15]))

	.dataa(gnd),
	.datab(\prif.rdat1_ex [15]),
	.datac(prifdmemaddr_15),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hF0CC;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N30
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (ptAScr & (!always02 & ((\Mux149~1_combout )))) # (!ptAScr & (((\Mux16~0_combout ))))

	.dataa(\HU|always0~6_combout ),
	.datab(\Mux16~0_combout ),
	.datac(\HU|ptAScr~4_combout ),
	.datad(\Mux149~1_combout ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'h5C0C;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N4
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (always02 & (prifdmemaddr_14)) # (!always02 & ((\prif.rdat1_ex [14])))

	.dataa(gnd),
	.datab(prifdmemaddr_14),
	.datac(\prif.rdat1_ex [14]),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hCCF0;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N18
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (ptAScr & (\Mux150~1_combout  & (!always02))) # (!ptAScr & (((\Mux17~0_combout ))))

	.dataa(\Mux150~1_combout ),
	.datab(\HU|always0~6_combout ),
	.datac(\Mux17~0_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'h22F0;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N4
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (always02 & (prifdmemaddr_13)) # (!always02 & ((\prif.rdat1_ex [13])))

	.dataa(prifdmemaddr_13),
	.datab(\prif.rdat1_ex [13]),
	.datac(gnd),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hAACC;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N30
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (ptAScr & (!always02 & (\Mux151~1_combout ))) # (!ptAScr & (((\Mux18~0_combout ))))

	.dataa(\HU|always0~6_combout ),
	.datab(\Mux151~1_combout ),
	.datac(\Mux18~0_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'h44F0;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N12
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (always02 & ((prifdmemaddr_11))) # (!always02 & (\prif.rdat1_ex [11]))

	.dataa(\HU|always0~6_combout ),
	.datab(gnd),
	.datac(\prif.rdat1_ex [11]),
	.datad(prifdmemaddr_11),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hFA50;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N14
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (ptAScr & (((\Mux153~1_combout  & !always02)))) # (!ptAScr & (\Mux20~0_combout ))

	.dataa(\Mux20~0_combout ),
	.datab(\Mux153~1_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'h0CAA;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N24
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (!always02 & (ptAScr & \Mux152~1_combout ))

	.dataa(gnd),
	.datab(\HU|always0~6_combout ),
	.datac(\HU|ptAScr~4_combout ),
	.datad(\Mux152~1_combout ),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'h3000;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N22
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (!ptAScr & ((always02 & (prifdmemaddr_12)) # (!always02 & ((\prif.rdat1_ex [12])))))

	.dataa(prifdmemaddr_12),
	.datab(\HU|ptAScr~4_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\prif.rdat1_ex [12]),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'h2320;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N10
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (always02 & (prifdmemaddr_10)) # (!always02 & ((\prif.rdat1_ex [10])))

	.dataa(\HU|always0~6_combout ),
	.datab(prifdmemaddr_10),
	.datac(gnd),
	.datad(\prif.rdat1_ex [10]),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hDD88;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N28
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (ptAScr & (((\Mux154~1_combout  & !always02)))) # (!ptAScr & (\Mux21~0_combout ))

	.dataa(\Mux21~0_combout ),
	.datab(\Mux154~1_combout ),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'h0CAA;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N14
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (always02 & ((prifdmemaddr_9))) # (!always02 & (\prif.rdat1_ex [9]))

	.dataa(\HU|always0~6_combout ),
	.datab(gnd),
	.datac(\prif.rdat1_ex [9]),
	.datad(prifdmemaddr_9),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hFA50;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N20
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (ptAScr & (!always02 & ((\Mux155~1_combout )))) # (!ptAScr & (((\Mux22~0_combout ))))

	.dataa(\HU|always0~6_combout ),
	.datab(\Mux22~0_combout ),
	.datac(\Mux155~1_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'h50CC;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N4
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (always02 & ((ptAScr & ((\prif.imm_mem [2]))) # (!ptAScr & (prifdmemaddr_18)))) # (!always02 & (((ptAScr))))

	.dataa(prifdmemaddr_18),
	.datab(\prif.imm_mem [2]),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hCFA0;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N26
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (always02 & (((\Mux13~0_combout )))) # (!always02 & ((\Mux13~0_combout  & ((\Mux146~1_combout ))) # (!\Mux13~0_combout  & (\prif.rdat1_ex [18]))))

	.dataa(\HU|always0~6_combout ),
	.datab(\prif.rdat1_ex [18]),
	.datac(\Mux13~0_combout ),
	.datad(\Mux146~1_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hF4A4;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N24
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (always02 & (((ptAScr)))) # (!always02 & ((ptAScr & (\Mux147~1_combout )) # (!ptAScr & ((\prif.rdat1_ex [17])))))

	.dataa(\Mux147~1_combout ),
	.datab(\prif.rdat1_ex [17]),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hFA0C;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N30
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (always02 & ((\Mux14~0_combout  & (\prif.imm_mem [1])) # (!\Mux14~0_combout  & ((prifdmemaddr_17))))) # (!always02 & (((\Mux14~0_combout ))))

	.dataa(\prif.imm_mem [1]),
	.datab(prifdmemaddr_17),
	.datac(\HU|always0~6_combout ),
	.datad(\Mux14~0_combout ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hAFC0;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N10
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (always02 & ((ptAScr) # ((prifdmemaddr_20)))) # (!always02 & (!ptAScr & ((\prif.rdat1_ex [20]))))

	.dataa(\HU|always0~6_combout ),
	.datab(\HU|ptAScr~4_combout ),
	.datac(prifdmemaddr_20),
	.datad(\prif.rdat1_ex [20]),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hB9A8;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N24
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (ptAScr & ((\Mux11~0_combout  & (\prif.imm_mem [4])) # (!\Mux11~0_combout  & ((\Mux144~1_combout ))))) # (!ptAScr & (((\Mux11~0_combout ))))

	.dataa(\prif.imm_mem [4]),
	.datab(\HU|ptAScr~4_combout ),
	.datac(\Mux144~1_combout ),
	.datad(\Mux11~0_combout ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hBBC0;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N24
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (ptAScr & ((\Mux145~1_combout ) # ((always02)))) # (!ptAScr & (((\prif.rdat1_ex [19] & !always02))))

	.dataa(\HU|ptAScr~4_combout ),
	.datab(\Mux145~1_combout ),
	.datac(\prif.rdat1_ex [19]),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hAAD8;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N30
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (always02 & ((\Mux12~0_combout  & ((\prif.imm_mem [3]))) # (!\Mux12~0_combout  & (prifdmemaddr_19)))) # (!always02 & (((\Mux12~0_combout ))))

	.dataa(\HU|always0~6_combout ),
	.datab(prifdmemaddr_19),
	.datac(\prif.imm_mem [3]),
	.datad(\Mux12~0_combout ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hF588;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N0
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (always02 & ((ptAScr) # ((prifdmemaddr_22)))) # (!always02 & (!ptAScr & ((\prif.rdat1_ex [22]))))

	.dataa(\HU|always0~6_combout ),
	.datab(\HU|ptAScr~4_combout ),
	.datac(prifdmemaddr_22),
	.datad(\prif.rdat1_ex [22]),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hB9A8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N26
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (ptAScr & ((\Mux9~0_combout  & ((\prif.imm_mem [6]))) # (!\Mux9~0_combout  & (\Mux142~1_combout )))) # (!ptAScr & (((\Mux9~0_combout ))))

	.dataa(\Mux142~1_combout ),
	.datab(\prif.imm_mem [6]),
	.datac(\HU|ptAScr~4_combout ),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hCFA0;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N30
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (ptAScr & (((\Mux143~1_combout ) # (always02)))) # (!ptAScr & (\prif.rdat1_ex [21] & ((!always02))))

	.dataa(\prif.rdat1_ex [21]),
	.datab(\Mux143~1_combout ),
	.datac(\HU|ptAScr~4_combout ),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hF0CA;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N16
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (\Mux10~0_combout  & ((\prif.imm_mem [5]) # ((!always02)))) # (!\Mux10~0_combout  & (((prifdmemaddr_21 & always02))))

	.dataa(\prif.imm_mem [5]),
	.datab(prifdmemaddr_21),
	.datac(\Mux10~0_combout ),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hACF0;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N4
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (always02 & ((prifdmemaddr_24) # ((ptAScr)))) # (!always02 & (((\prif.rdat1_ex [24] & !ptAScr))))

	.dataa(prifdmemaddr_24),
	.datab(\HU|always0~6_combout ),
	.datac(\prif.rdat1_ex [24]),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hCCB8;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N10
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (\Mux7~0_combout  & ((\prif.imm_mem [8]) # ((!ptAScr)))) # (!\Mux7~0_combout  & (((\Mux140~1_combout  & ptAScr))))

	.dataa(\prif.imm_mem [8]),
	.datab(\Mux140~1_combout ),
	.datac(\Mux7~0_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hACF0;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N16
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (ptAScr & ((\Mux141~1_combout ) # ((always02)))) # (!ptAScr & (((\prif.rdat1_ex [23] & !always02))))

	.dataa(\Mux141~1_combout ),
	.datab(\HU|ptAScr~4_combout ),
	.datac(\prif.rdat1_ex [23]),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hCCB8;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N6
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (always02 & ((\Mux8~0_combout  & (\prif.imm_mem [7])) # (!\Mux8~0_combout  & ((prifdmemaddr_23))))) # (!always02 & (((\Mux8~0_combout ))))

	.dataa(\HU|always0~6_combout ),
	.datab(\prif.imm_mem [7]),
	.datac(prifdmemaddr_23),
	.datad(\Mux8~0_combout ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hDDA0;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N24
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (always02 & (((ptAScr)))) # (!always02 & ((ptAScr & (\Mux133~1_combout )) # (!ptAScr & ((\prif.rdat1_ex [31])))))

	.dataa(\Mux133~1_combout ),
	.datab(\HU|always0~6_combout ),
	.datac(\prif.rdat1_ex [31]),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hEE30;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N18
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (always02 & ((\Mux0~0_combout  & ((\prif.imm_mem [15]))) # (!\Mux0~0_combout  & (prifdmemaddr_31)))) # (!always02 & (((\Mux0~0_combout ))))

	.dataa(prifdmemaddr_31),
	.datab(\prif.imm_mem [15]),
	.datac(\HU|always0~6_combout ),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hCFA0;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N6
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (always02 & (((prifdmemaddr_30) # (ptAScr)))) # (!always02 & (\prif.rdat1_ex [30] & ((!ptAScr))))

	.dataa(\prif.rdat1_ex [30]),
	.datab(prifdmemaddr_30),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hF0CA;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N12
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (ptAScr & ((\Mux1~0_combout  & ((\prif.imm_mem [14]))) # (!\Mux1~0_combout  & (\Mux134~1_combout )))) # (!ptAScr & (((\Mux1~0_combout ))))

	.dataa(\HU|ptAScr~4_combout ),
	.datab(\Mux134~1_combout ),
	.datac(\prif.imm_mem [14]),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hF588;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N18
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (always02 & (((ptAScr)))) # (!always02 & ((ptAScr & ((\Mux135~1_combout ))) # (!ptAScr & (\prif.rdat1_ex [29]))))

	.dataa(\HU|always0~6_combout ),
	.datab(\prif.rdat1_ex [29]),
	.datac(\HU|ptAScr~4_combout ),
	.datad(\Mux135~1_combout ),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hF4A4;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N4
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (always02 & ((\Mux2~0_combout  & (\prif.imm_mem [13])) # (!\Mux2~0_combout  & ((prifdmemaddr_29))))) # (!always02 & (((\Mux2~0_combout ))))

	.dataa(\HU|always0~6_combout ),
	.datab(\prif.imm_mem [13]),
	.datac(prifdmemaddr_29),
	.datad(\Mux2~0_combout ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hDDA0;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N4
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (always02 & ((prifdmemaddr_26) # ((ptAScr)))) # (!always02 & (((!ptAScr & \prif.rdat1_ex [26]))))

	.dataa(prifdmemaddr_26),
	.datab(\HU|always0~6_combout ),
	.datac(\HU|ptAScr~4_combout ),
	.datad(\prif.rdat1_ex [26]),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hCBC8;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N18
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (ptAScr & ((\Mux5~0_combout  & (\prif.imm_mem [10])) # (!\Mux5~0_combout  & ((\Mux138~1_combout ))))) # (!ptAScr & (((\Mux5~0_combout ))))

	.dataa(\prif.imm_mem [10]),
	.datab(\HU|ptAScr~4_combout ),
	.datac(\Mux5~0_combout ),
	.datad(\Mux138~1_combout ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hBCB0;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N18
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (always02 & (((ptAScr)))) # (!always02 & ((ptAScr & (\Mux139~1_combout )) # (!ptAScr & ((\prif.rdat1_ex [25])))))

	.dataa(\Mux139~1_combout ),
	.datab(\prif.rdat1_ex [25]),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hFA0C;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N28
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (always02 & ((\Mux6~0_combout  & (\prif.imm_mem [9])) # (!\Mux6~0_combout  & ((prifdmemaddr_25))))) # (!always02 & (((\Mux6~0_combout ))))

	.dataa(\HU|always0~6_combout ),
	.datab(\prif.imm_mem [9]),
	.datac(prifdmemaddr_25),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hDDA0;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N6
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (always02 & (((prifdmemaddr_28) # (ptAScr)))) # (!always02 & (\prif.rdat1_ex [28] & ((!ptAScr))))

	.dataa(\prif.rdat1_ex [28]),
	.datab(prifdmemaddr_28),
	.datac(\HU|always0~6_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hF0CA;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N24
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (\Mux3~0_combout  & (((\prif.imm_mem [12]) # (!ptAScr)))) # (!\Mux3~0_combout  & (\Mux136~1_combout  & ((ptAScr))))

	.dataa(\Mux3~0_combout ),
	.datab(\Mux136~1_combout ),
	.datac(\prif.imm_mem [12]),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hE4AA;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N30
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (always02 & (((ptAScr)))) # (!always02 & ((ptAScr & ((\Mux137~1_combout ))) # (!ptAScr & (\prif.rdat1_ex [27]))))

	.dataa(\prif.rdat1_ex [27]),
	.datab(\HU|always0~6_combout ),
	.datac(\Mux137~1_combout ),
	.datad(\HU|ptAScr~4_combout ),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hFC22;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N8
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (\Mux4~0_combout  & ((\prif.imm_mem [11]) # ((!always02)))) # (!\Mux4~0_combout  & (((prifdmemaddr_27 & always02))))

	.dataa(\prif.imm_mem [11]),
	.datab(prifdmemaddr_27),
	.datac(\Mux4~0_combout ),
	.datad(\HU|always0~6_combout ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hACF0;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y24_N13
dffeas \prif.ALUOP_ex[0] (
	.clk(CLK),
	.d(\PR|ALUOP_ex~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.ALUOP_ex [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.ALUOP_ex[0] .is_wysiwyg = "true";
defparam \prif.ALUOP_ex[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N4
cycloneive_lcell_comb \Equal1~0 (
// Equation(s):
// \Equal1~0_combout  = (!\prif.opcode_mem [3] & (!\prif.opcode_mem [4] & (!\prif.opcode_mem [5] & !\prif.opcode_mem [0])))

	.dataa(\prif.opcode_mem [3]),
	.datab(\prif.opcode_mem [4]),
	.datac(\prif.opcode_mem [5]),
	.datad(\prif.opcode_mem [0]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0001;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N8
cycloneive_lcell_comb \Equal1~1 (
// Equation(s):
// \Equal1~1_combout  = (!\prif.opcode_mem [1] & (\Equal1~0_combout  & \prif.opcode_mem [2]))

	.dataa(gnd),
	.datab(\prif.opcode_mem [1]),
	.datac(\Equal1~0_combout ),
	.datad(\prif.opcode_mem [2]),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'h3000;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N16
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (always02 & (prifdmemaddr_12)) # (!always02 & ((\prif.rdat1_ex [12])))

	.dataa(prifdmemaddr_12),
	.datab(gnd),
	.datac(\HU|always0~6_combout ),
	.datad(\prif.rdat1_ex [12]),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hAFA0;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N26
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (ptAScr & (\Mux152~1_combout  & (!always02))) # (!ptAScr & (((\Mux19~2_combout ))))

	.dataa(\Mux152~1_combout ),
	.datab(\HU|always0~6_combout ),
	.datac(\HU|ptAScr~4_combout ),
	.datad(\Mux19~2_combout ),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'h2F20;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y28_N29
dffeas \prif.pc_mem[1] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[1]~4_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[1] .is_wysiwyg = "true";
defparam \prif.pc_mem[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N30
cycloneive_lcell_comb \prif.rs_ex[0]~0 (
// Equation(s):
// \prif.rs_ex[0]~0_combout  = ((ccifiwait_0) # (flush_idex)) # (!\nRST~input_o )

	.dataa(nRST),
	.datab(gnd),
	.datac(ccifiwait_0),
	.datad(\HU|flush_idex~0_combout ),
	.cin(gnd),
	.combout(\prif.rs_ex[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \prif.rs_ex[0]~0 .lut_mask = 16'hFFF5;
defparam \prif.rs_ex[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X53_Y28_N27
dffeas \prif.pc_mem[0] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[0]~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[0] .is_wysiwyg = "true";
defparam \prif.pc_mem[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y34_N9
dffeas \prif.pc_mem[3] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[3]~6_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[3] .is_wysiwyg = "true";
defparam \prif.pc_mem[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N27
dffeas \prif.pc_mem[2] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[2]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[2] .is_wysiwyg = "true";
defparam \prif.pc_mem[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y27_N25
dffeas \prif.pc_mem[4] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[4]~8_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[4] .is_wysiwyg = "true";
defparam \prif.pc_mem[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N11
dffeas \prif.pc_mem[5] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[5]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[5] .is_wysiwyg = "true";
defparam \prif.pc_mem[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N27
dffeas \prif.pc_mem[15] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[15]~10_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[15] .is_wysiwyg = "true";
defparam \prif.pc_mem[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y34_N19
dffeas \prif.pc_mem[14] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[14]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[14] .is_wysiwyg = "true";
defparam \prif.pc_mem[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N9
dffeas \prif.pc_mem[13] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[13]~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[13] .is_wysiwyg = "true";
defparam \prif.pc_mem[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N17
dffeas \prif.pc_mem[12] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[12]~13_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[12] .is_wysiwyg = "true";
defparam \prif.pc_mem[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N15
dffeas \prif.pc_mem[11] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[11]~14_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[11] .is_wysiwyg = "true";
defparam \prif.pc_mem[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N25
dffeas \prif.pc_mem[10] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[10]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[10] .is_wysiwyg = "true";
defparam \prif.pc_mem[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N1
dffeas \prif.pc_mem[9] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[9]~16_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[9] .is_wysiwyg = "true";
defparam \prif.pc_mem[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N3
dffeas \prif.pc_mem[6] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[6]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[6] .is_wysiwyg = "true";
defparam \prif.pc_mem[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N21
dffeas \prif.pc_mem[27] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[27]~18_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[27] .is_wysiwyg = "true";
defparam \prif.pc_mem[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N19
dffeas \prif.pc_mem[23] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[23]~19_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[23] .is_wysiwyg = "true";
defparam \prif.pc_mem[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N17
dffeas \prif.pc_mem[18] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[18]~20_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[18] .is_wysiwyg = "true";
defparam \prif.pc_mem[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N31
dffeas \prif.pc_mem[24] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[24]~21_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[24] .is_wysiwyg = "true";
defparam \prif.pc_mem[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y27_N21
dffeas \prif.pc_mem[16] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[16]~22_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[16] .is_wysiwyg = "true";
defparam \prif.pc_mem[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N9
dffeas \prif.pc_mem[19] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[19]~23_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[19] .is_wysiwyg = "true";
defparam \prif.pc_mem[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N23
dffeas \prif.pc_mem[17] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[17]~24_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[17] .is_wysiwyg = "true";
defparam \prif.pc_mem[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N5
dffeas \prif.pc_mem[21] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[21]~25_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[21] .is_wysiwyg = "true";
defparam \prif.pc_mem[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N15
dffeas \prif.pc_mem[20] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[20]~26_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[20] .is_wysiwyg = "true";
defparam \prif.pc_mem[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y32_N7
dffeas \prif.pc_mem[26] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[26]~27_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[26] .is_wysiwyg = "true";
defparam \prif.pc_mem[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N21
dffeas \prif.pc_mem[8] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[8]~28_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[8] .is_wysiwyg = "true";
defparam \prif.pc_mem[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y33_N7
dffeas \prif.pc_mem[7] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[7]~29_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[7] .is_wysiwyg = "true";
defparam \prif.pc_mem[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y31_N23
dffeas \prif.pc_mem[22] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[22]~30_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[22] .is_wysiwyg = "true";
defparam \prif.pc_mem[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y33_N3
dffeas \prif.pc_mem[25] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[25]~31_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[25] .is_wysiwyg = "true";
defparam \prif.pc_mem[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N20
cycloneive_lcell_comb \prif.pc_mem[15]~0 (
// Equation(s):
// \prif.pc_mem[15]~0_combout  = (((always1) # (always01)) # (!always1)) # (!\nRST~input_o )

	.dataa(nRST),
	.datab(always1),
	.datac(\HU|always1~5_combout ),
	.datad(always01),
	.cin(gnd),
	.combout(\prif.pc_mem[15]~0_combout ),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[15]~0 .lut_mask = 16'hFFF7;
defparam \prif.pc_mem[15]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N10
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (\Mux60~0_combout ) # ((prifdmemaddr_3 & (!always01 & ptBScr)))

	.dataa(prifdmemaddr_3),
	.datab(\HU|always0~5_combout ),
	.datac(\Mux60~0_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hF2F0;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N4
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (\Mux59~0_combout ) # ((ptBScr & (prifdmemaddr_4 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_4),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux59~0_combout ),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hFF08;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N20
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (\Mux58~0_combout ) # ((!always01 & (ptBScr & prifdmemaddr_5)))

	.dataa(\Mux58~0_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(\HU|ptBScr~1_combout ),
	.datad(prifdmemaddr_5),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hBAAA;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N24
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (\Mux57~0_combout ) # ((ptBScr & (prifdmemaddr_6 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_6),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux57~0_combout ),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hFF08;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N22
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (\Mux56~0_combout ) # ((ptBScr & (prifdmemaddr_7 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_7),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux56~0_combout ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hFF08;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N0
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (\Mux55~0_combout ) # ((!always01 & (ptBScr & prifdmemaddr_8)))

	.dataa(\Mux55~0_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(\HU|ptBScr~1_combout ),
	.datad(prifdmemaddr_8),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hBAAA;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N14
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (\Mux54~0_combout ) # ((prifdmemaddr_9 & (!always01 & ptBScr)))

	.dataa(prifdmemaddr_9),
	.datab(\HU|always0~5_combout ),
	.datac(\HU|ptBScr~1_combout ),
	.datad(\Mux54~0_combout ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hFF20;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N6
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (\Mux53~0_combout ) # ((ptBScr & (!always01 & prifdmemaddr_10)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(\HU|always0~5_combout ),
	.datac(\Mux53~0_combout ),
	.datad(prifdmemaddr_10),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hF2F0;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N10
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (\Mux52~0_combout ) # ((prifdmemaddr_11 & (!always01 & ptBScr)))

	.dataa(prifdmemaddr_11),
	.datab(\Mux52~0_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hCECC;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N12
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (\Mux51~0_combout ) # ((ptBScr & (prifdmemaddr_12 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_12),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux51~0_combout ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hFF08;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N8
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (\Mux50~0_combout ) # ((!always01 & (ptBScr & prifdmemaddr_13)))

	.dataa(\HU|always0~5_combout ),
	.datab(\HU|ptBScr~1_combout ),
	.datac(prifdmemaddr_13),
	.datad(\Mux50~0_combout ),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hFF40;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N20
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (\Mux49~0_combout ) # ((ptBScr & (prifdmemaddr_14 & !always01)))

	.dataa(\HU|ptBScr~1_combout ),
	.datab(prifdmemaddr_14),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux49~0_combout ),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hFF08;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N10
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (ptBScr & ((prifdmemaddr_15))) # (!ptBScr & (\prif.rdat2_ex [15]))

	.dataa(\prif.rdat2_ex [15]),
	.datab(gnd),
	.datac(prifdmemaddr_15),
	.datad(\HU|ptBScr~1_combout ),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hF0AA;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N20
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (always01 & (((!ptBScr & \Mux149~1_combout )))) # (!always01 & (\Mux48~0_combout ))

	.dataa(\Mux48~0_combout ),
	.datab(\HU|ptBScr~1_combout ),
	.datac(\HU|always0~5_combout ),
	.datad(\Mux149~1_combout ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'h3A0A;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y29_N3
dffeas \prif.halt_wb (
	.clk(CLK),
	.d(\PR|halt_wb~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.halt_wb~q ),
	.prn(vcc));
// synopsys translate_off
defparam \prif.halt_wb .is_wysiwyg = "true";
defparam \prif.halt_wb .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N26
cycloneive_lcell_comb \Mux90~3 (
// Equation(s):
// \Mux90~3_combout  = (\prif.ALUScr_ex [0] & (\prif.imm_ex [5])) # (!\prif.ALUScr_ex [0] & (((!\prif.ALUScr_ex [1] & \Mux90~2_combout ))))

	.dataa(\prif.imm_ex [5]),
	.datab(\prif.ALUScr_ex [1]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux90~2_combout ),
	.cin(gnd),
	.combout(\Mux90~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux90~3 .lut_mask = 16'hA3A0;
defparam \Mux90~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N6
cycloneive_lcell_comb \Mux80~4 (
// Equation(s):
// \Mux80~4_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [15])))) # (!\prif.ALUScr_ex [0] & (!\prif.ALUScr_ex [1] & ((\Mux80~3_combout ))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.imm_ex [15]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux80~3_combout ),
	.cin(gnd),
	.combout(\Mux80~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux80~4 .lut_mask = 16'hC5C0;
defparam \Mux80~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N6
cycloneive_lcell_comb \Mux81~3 (
// Equation(s):
// \Mux81~3_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [14])))) # (!\prif.ALUScr_ex [0] & (!\prif.ALUScr_ex [1] & ((\Mux81~2_combout ))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.ALUScr_ex [0]),
	.datac(\prif.imm_ex [14]),
	.datad(\Mux81~2_combout ),
	.cin(gnd),
	.combout(\Mux81~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux81~3 .lut_mask = 16'hD1C0;
defparam \Mux81~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N6
cycloneive_lcell_comb \Mux82~3 (
// Equation(s):
// \Mux82~3_combout  = (\prif.ALUScr_ex [0] & (\prif.imm_ex [13])) # (!\prif.ALUScr_ex [0] & (((!\prif.ALUScr_ex [1] & \Mux82~2_combout ))))

	.dataa(\prif.imm_ex [13]),
	.datab(\prif.ALUScr_ex [1]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux82~2_combout ),
	.cin(gnd),
	.combout(\Mux82~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux82~3 .lut_mask = 16'hA3A0;
defparam \Mux82~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N18
cycloneive_lcell_comb \Mux83~3 (
// Equation(s):
// \Mux83~3_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [12])))) # (!\prif.ALUScr_ex [0] & (!\prif.ALUScr_ex [1] & ((\Mux83~2_combout ))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.imm_ex [12]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux83~2_combout ),
	.cin(gnd),
	.combout(\Mux83~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux83~3 .lut_mask = 16'hC5C0;
defparam \Mux83~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N14
cycloneive_lcell_comb \Mux84~3 (
// Equation(s):
// \Mux84~3_combout  = (\prif.ALUScr_ex [0] & (\prif.imm_ex [11])) # (!\prif.ALUScr_ex [0] & (((!\prif.ALUScr_ex [1] & \Mux84~2_combout ))))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.imm_ex [11]),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\Mux84~2_combout ),
	.cin(gnd),
	.combout(\Mux84~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux84~3 .lut_mask = 16'h8D88;
defparam \Mux84~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N4
cycloneive_lcell_comb \Mux85~3 (
// Equation(s):
// \Mux85~3_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [10])))) # (!\prif.ALUScr_ex [0] & (!\prif.ALUScr_ex [1] & ((\Mux85~2_combout ))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.imm_ex [10]),
	.datac(\prif.ALUScr_ex [0]),
	.datad(\Mux85~2_combout ),
	.cin(gnd),
	.combout(\Mux85~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux85~3 .lut_mask = 16'hC5C0;
defparam \Mux85~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N10
cycloneive_lcell_comb \Mux86~3 (
// Equation(s):
// \Mux86~3_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [9])))) # (!\prif.ALUScr_ex [0] & (\Mux86~2_combout  & ((!\prif.ALUScr_ex [1]))))

	.dataa(\Mux86~2_combout ),
	.datab(\prif.ALUScr_ex [0]),
	.datac(\prif.imm_ex [9]),
	.datad(\prif.ALUScr_ex [1]),
	.cin(gnd),
	.combout(\Mux86~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux86~3 .lut_mask = 16'hC0E2;
defparam \Mux86~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N6
cycloneive_lcell_comb \Mux89~4 (
// Equation(s):
// \Mux89~4_combout  = (\prif.ALUScr_ex [0] & (\prif.imm_ex [6])) # (!\prif.ALUScr_ex [0] & (((!\prif.ALUScr_ex [1] & \Mux89~3_combout ))))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.imm_ex [6]),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\Mux89~3_combout ),
	.cin(gnd),
	.combout(\Mux89~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux89~4 .lut_mask = 16'h8D88;
defparam \Mux89~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N28
cycloneive_lcell_comb \Mux87~3 (
// Equation(s):
// \Mux87~3_combout  = (\prif.ALUScr_ex [0] & (\prif.imm_ex [8])) # (!\prif.ALUScr_ex [0] & (((!\prif.ALUScr_ex [1] & \Mux87~2_combout ))))

	.dataa(\prif.ALUScr_ex [0]),
	.datab(\prif.imm_ex [8]),
	.datac(\prif.ALUScr_ex [1]),
	.datad(\Mux87~2_combout ),
	.cin(gnd),
	.combout(\Mux87~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux87~3 .lut_mask = 16'h8D88;
defparam \Mux87~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N10
cycloneive_lcell_comb \Mux88~3 (
// Equation(s):
// \Mux88~3_combout  = (\prif.ALUScr_ex [0] & (((\prif.imm_ex [7])))) # (!\prif.ALUScr_ex [0] & (!\prif.ALUScr_ex [1] & ((\Mux88~2_combout ))))

	.dataa(\prif.ALUScr_ex [1]),
	.datab(\prif.imm_ex [7]),
	.datac(\Mux88~2_combout ),
	.datad(\prif.ALUScr_ex [0]),
	.cin(gnd),
	.combout(\Mux88~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux88~3 .lut_mask = 16'hCC50;
defparam \Mux88~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N4
cycloneive_lcell_comb \prif.ALUScr_ex[0]~feeder (
// Equation(s):
// \prif.ALUScr_ex[0]~feeder_combout  = ALUScr_ex1

	.dataa(\PR|ALUScr_ex~12_combout ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\prif.ALUScr_ex[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \prif.ALUScr_ex[0]~feeder .lut_mask = 16'hAAAA;
defparam \prif.ALUScr_ex[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y25_N25
dffeas \prif.dmemaddr[1] (
	.clk(CLK),
	.d(\PR|dmemaddr~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_1),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[1] .is_wysiwyg = "true";
defparam \prif.dmemaddr[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N17
dffeas \pc[1] (
	.clk(CLK),
	.d(\Mux131~0_combout ),
	.asdata(\prif.pc_bran_mem [1]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\prif.PCScr_mem [1]),
	.ena(\pc[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_1),
	.prn(vcc));
// synopsys translate_off
defparam \pc[1] .is_wysiwyg = "true";
defparam \pc[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y29_N29
dffeas \prif.dmemren (
	.clk(CLK),
	.d(\PR|dmemren~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemren),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemren .is_wysiwyg = "true";
defparam \prif.dmemren .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y29_N15
dffeas \prif.dmemwen (
	.clk(CLK),
	.d(\PR|dmemwen~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemwen),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemwen .is_wysiwyg = "true";
defparam \prif.dmemwen .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y25_N5
dffeas \prif.dmemaddr[0] (
	.clk(CLK),
	.d(\PR|dmemaddr~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_0),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[0] .is_wysiwyg = "true";
defparam \prif.dmemaddr[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N31
dffeas \pc[0] (
	.clk(CLK),
	.d(\Mux132~0_combout ),
	.asdata(\prif.pc_bran_mem [0]),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(!\prif.PCScr_mem [1]),
	.ena(\pc[1]~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_0),
	.prn(vcc));
// synopsys translate_off
defparam \pc[0] .is_wysiwyg = "true";
defparam \pc[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y25_N31
dffeas \prif.dmemaddr[3] (
	.clk(CLK),
	.d(\PR|dmemaddr~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_3),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[3] .is_wysiwyg = "true";
defparam \prif.dmemaddr[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y25_N1
dffeas \prif.dmemaddr[2] (
	.clk(CLK),
	.d(\PR|dmemaddr~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_2),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[2] .is_wysiwyg = "true";
defparam \prif.dmemaddr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N17
dffeas \prif.dmemaddr[5] (
	.clk(CLK),
	.d(\PR|dmemaddr~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_5),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[5] .is_wysiwyg = "true";
defparam \prif.dmemaddr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N19
dffeas \prif.dmemaddr[4] (
	.clk(CLK),
	.d(\PR|dmemaddr~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_4),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[4] .is_wysiwyg = "true";
defparam \prif.dmemaddr[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N5
dffeas \prif.dmemaddr[7] (
	.clk(CLK),
	.d(\PR|dmemaddr~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_7),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[7] .is_wysiwyg = "true";
defparam \prif.dmemaddr[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N15
dffeas \prif.dmemaddr[6] (
	.clk(CLK),
	.d(\PR|dmemaddr~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_6),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[6] .is_wysiwyg = "true";
defparam \prif.dmemaddr[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N9
dffeas \prif.dmemaddr[9] (
	.clk(CLK),
	.d(\PR|dmemaddr~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_9),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[9] .is_wysiwyg = "true";
defparam \prif.dmemaddr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N23
dffeas \prif.dmemaddr[8] (
	.clk(CLK),
	.d(\PR|dmemaddr~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_8),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[8] .is_wysiwyg = "true";
defparam \prif.dmemaddr[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y25_N23
dffeas \prif.dmemaddr[11] (
	.clk(CLK),
	.d(\PR|dmemaddr~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_11),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[11] .is_wysiwyg = "true";
defparam \prif.dmemaddr[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y25_N17
dffeas \prif.dmemaddr[10] (
	.clk(CLK),
	.d(\PR|dmemaddr~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_10),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[10] .is_wysiwyg = "true";
defparam \prif.dmemaddr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N13
dffeas \prif.dmemaddr[13] (
	.clk(CLK),
	.d(\PR|dmemaddr~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_13),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[13] .is_wysiwyg = "true";
defparam \prif.dmemaddr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N31
dffeas \prif.dmemaddr[12] (
	.clk(CLK),
	.d(\PR|dmemaddr~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_12),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[12] .is_wysiwyg = "true";
defparam \prif.dmemaddr[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y26_N9
dffeas \prif.dmemaddr[15] (
	.clk(CLK),
	.d(\PR|dmemaddr~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_15),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[15] .is_wysiwyg = "true";
defparam \prif.dmemaddr[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y26_N9
dffeas \prif.dmemaddr[14] (
	.clk(CLK),
	.d(\PR|dmemaddr~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_14),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[14] .is_wysiwyg = "true";
defparam \prif.dmemaddr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N5
dffeas \prif.dmemaddr[23] (
	.clk(CLK),
	.d(\PR|dmemaddr~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_23),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[23] .is_wysiwyg = "true";
defparam \prif.dmemaddr[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N15
dffeas \prif.dmemaddr[22] (
	.clk(CLK),
	.d(\PR|dmemaddr~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_22),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[22] .is_wysiwyg = "true";
defparam \prif.dmemaddr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N29
dffeas \prif.dmemaddr[21] (
	.clk(CLK),
	.d(\PR|dmemaddr~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_21),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[21] .is_wysiwyg = "true";
defparam \prif.dmemaddr[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y31_N9
dffeas \prif.dmemaddr[29] (
	.clk(CLK),
	.d(\PR|dmemaddr~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_29),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[29] .is_wysiwyg = "true";
defparam \prif.dmemaddr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y25_N27
dffeas \prif.dmemaddr[28] (
	.clk(CLK),
	.d(\PR|dmemaddr~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_28),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[28] .is_wysiwyg = "true";
defparam \prif.dmemaddr[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y28_N9
dffeas \prif.dmemaddr[31] (
	.clk(CLK),
	.d(\PR|dmemaddr~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_31),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[31] .is_wysiwyg = "true";
defparam \prif.dmemaddr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N1
dffeas \prif.dmemaddr[30] (
	.clk(CLK),
	.d(\PR|dmemaddr~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_30),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[30] .is_wysiwyg = "true";
defparam \prif.dmemaddr[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N1
dffeas \prif.dmemaddr[20] (
	.clk(CLK),
	.d(\PR|dmemaddr~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_20),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[20] .is_wysiwyg = "true";
defparam \prif.dmemaddr[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N11
dffeas \prif.dmemaddr[17] (
	.clk(CLK),
	.d(\PR|dmemaddr~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_17),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[17] .is_wysiwyg = "true";
defparam \prif.dmemaddr[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N13
dffeas \prif.dmemaddr[16] (
	.clk(CLK),
	.d(\PR|dmemaddr~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_16),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[16] .is_wysiwyg = "true";
defparam \prif.dmemaddr[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N1
dffeas \prif.dmemaddr[19] (
	.clk(CLK),
	.d(\PR|dmemaddr~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_19),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[19] .is_wysiwyg = "true";
defparam \prif.dmemaddr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y25_N5
dffeas \prif.dmemaddr[18] (
	.clk(CLK),
	.d(\PR|dmemaddr~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_18),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[18] .is_wysiwyg = "true";
defparam \prif.dmemaddr[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N17
dffeas \prif.dmemaddr[25] (
	.clk(CLK),
	.d(\PR|dmemaddr~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_25),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[25] .is_wysiwyg = "true";
defparam \prif.dmemaddr[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y25_N13
dffeas \prif.dmemaddr[24] (
	.clk(CLK),
	.d(\PR|dmemaddr~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_24),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[24] .is_wysiwyg = "true";
defparam \prif.dmemaddr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y26_N29
dffeas \prif.dmemaddr[27] (
	.clk(CLK),
	.d(\PR|dmemaddr~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_27),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[27] .is_wysiwyg = "true";
defparam \prif.dmemaddr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N13
dffeas \prif.dmemaddr[26] (
	.clk(CLK),
	.d(\PR|dmemaddr~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemaddr_26),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemaddr[26] .is_wysiwyg = "true";
defparam \prif.dmemaddr[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y29_N11
dffeas \prif.dmemstore[0] (
	.clk(CLK),
	.d(\PR|dmemstore~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_0),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[0] .is_wysiwyg = "true";
defparam \prif.dmemstore[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y26_N19
dffeas \prif.dmemstore[1] (
	.clk(CLK),
	.d(\PR|dmemstore~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_1),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[1] .is_wysiwyg = "true";
defparam \prif.dmemstore[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y26_N21
dffeas \prif.dmemstore[2] (
	.clk(CLK),
	.d(\PR|dmemstore~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_2),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[2] .is_wysiwyg = "true";
defparam \prif.dmemstore[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y26_N27
dffeas \prif.dmemstore[3] (
	.clk(CLK),
	.d(\PR|dmemstore~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_3),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[3] .is_wysiwyg = "true";
defparam \prif.dmemstore[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y26_N17
dffeas \prif.dmemstore[4] (
	.clk(CLK),
	.d(\PR|dmemstore~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_4),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[4] .is_wysiwyg = "true";
defparam \prif.dmemstore[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y26_N3
dffeas \prif.dmemstore[5] (
	.clk(CLK),
	.d(\PR|dmemstore~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_5),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[5] .is_wysiwyg = "true";
defparam \prif.dmemstore[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y26_N25
dffeas \prif.dmemstore[6] (
	.clk(CLK),
	.d(\PR|dmemstore~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_6),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[6] .is_wysiwyg = "true";
defparam \prif.dmemstore[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y29_N21
dffeas \prif.dmemstore[7] (
	.clk(CLK),
	.d(\PR|dmemstore~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_7),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[7] .is_wysiwyg = "true";
defparam \prif.dmemstore[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y26_N11
dffeas \prif.dmemstore[8] (
	.clk(CLK),
	.d(\PR|dmemstore~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_8),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[8] .is_wysiwyg = "true";
defparam \prif.dmemstore[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y29_N19
dffeas \prif.dmemstore[9] (
	.clk(CLK),
	.d(\PR|dmemstore~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_9),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[9] .is_wysiwyg = "true";
defparam \prif.dmemstore[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N21
dffeas \prif.dmemstore[10] (
	.clk(CLK),
	.d(\PR|dmemstore~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_10),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[10] .is_wysiwyg = "true";
defparam \prif.dmemstore[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N7
dffeas \prif.dmemstore[11] (
	.clk(CLK),
	.d(\PR|dmemstore~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_11),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[11] .is_wysiwyg = "true";
defparam \prif.dmemstore[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N29
dffeas \prif.dmemstore[12] (
	.clk(CLK),
	.d(\PR|dmemstore~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_12),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[12] .is_wysiwyg = "true";
defparam \prif.dmemstore[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y26_N13
dffeas \prif.dmemstore[13] (
	.clk(CLK),
	.d(\PR|dmemstore~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_13),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[13] .is_wysiwyg = "true";
defparam \prif.dmemstore[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N19
dffeas \prif.dmemstore[14] (
	.clk(CLK),
	.d(\PR|dmemstore~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_14),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[14] .is_wysiwyg = "true";
defparam \prif.dmemstore[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N25
dffeas \prif.dmemstore[15] (
	.clk(CLK),
	.d(\PR|dmemstore~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_15),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[15] .is_wysiwyg = "true";
defparam \prif.dmemstore[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N11
dffeas \prif.dmemstore[16] (
	.clk(CLK),
	.d(\PR|dmemstore~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_16),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[16] .is_wysiwyg = "true";
defparam \prif.dmemstore[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N13
dffeas \prif.dmemstore[17] (
	.clk(CLK),
	.d(\PR|dmemstore~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_17),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[17] .is_wysiwyg = "true";
defparam \prif.dmemstore[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y30_N3
dffeas \prif.dmemstore[18] (
	.clk(CLK),
	.d(\PR|dmemstore~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_18),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[18] .is_wysiwyg = "true";
defparam \prif.dmemstore[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N21
dffeas \prif.dmemstore[19] (
	.clk(CLK),
	.d(\PR|dmemstore~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_19),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[19] .is_wysiwyg = "true";
defparam \prif.dmemstore[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N7
dffeas \prif.dmemstore[20] (
	.clk(CLK),
	.d(\PR|dmemstore~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_20),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[20] .is_wysiwyg = "true";
defparam \prif.dmemstore[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N13
dffeas \prif.dmemstore[21] (
	.clk(CLK),
	.d(\PR|dmemstore~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_21),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[21] .is_wysiwyg = "true";
defparam \prif.dmemstore[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N31
dffeas \prif.dmemstore[22] (
	.clk(CLK),
	.d(\PR|dmemstore~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_22),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[22] .is_wysiwyg = "true";
defparam \prif.dmemstore[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N11
dffeas \prif.dmemstore[23] (
	.clk(CLK),
	.d(\PR|dmemstore~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_23),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[23] .is_wysiwyg = "true";
defparam \prif.dmemstore[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y27_N1
dffeas \prif.dmemstore[24] (
	.clk(CLK),
	.d(\PR|dmemstore~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_24),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[24] .is_wysiwyg = "true";
defparam \prif.dmemstore[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N17
dffeas \prif.dmemstore[25] (
	.clk(CLK),
	.d(\PR|dmemstore~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_25),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[25] .is_wysiwyg = "true";
defparam \prif.dmemstore[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y27_N3
dffeas \prif.dmemstore[26] (
	.clk(CLK),
	.d(\PR|dmemstore~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_26),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[26] .is_wysiwyg = "true";
defparam \prif.dmemstore[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y26_N27
dffeas \prif.dmemstore[27] (
	.clk(CLK),
	.d(\PR|dmemstore~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_27),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[27] .is_wysiwyg = "true";
defparam \prif.dmemstore[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y26_N19
dffeas \prif.dmemstore[28] (
	.clk(CLK),
	.d(\PR|dmemstore~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_28),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[28] .is_wysiwyg = "true";
defparam \prif.dmemstore[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y30_N3
dffeas \prif.dmemstore[29] (
	.clk(CLK),
	.d(\PR|dmemstore~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_29),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[29] .is_wysiwyg = "true";
defparam \prif.dmemstore[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y28_N23
dffeas \prif.dmemstore[30] (
	.clk(CLK),
	.d(\PR|dmemstore~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_30),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[30] .is_wysiwyg = "true";
defparam \prif.dmemstore[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y29_N9
dffeas \prif.dmemstore[31] (
	.clk(CLK),
	.d(\PR|dmemstore~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(prifdmemstore_31),
	.prn(vcc));
// synopsys translate_off
defparam \prif.dmemstore[31] .is_wysiwyg = "true";
defparam \prif.dmemstore[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N1
dffeas \pc[3] (
	.clk(CLK),
	.d(\Mux129~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_3),
	.prn(vcc));
// synopsys translate_off
defparam \pc[3] .is_wysiwyg = "true";
defparam \pc[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N9
dffeas \pc[2] (
	.clk(CLK),
	.d(\Mux130~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_2),
	.prn(vcc));
// synopsys translate_off
defparam \pc[2] .is_wysiwyg = "true";
defparam \pc[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y28_N23
dffeas \pc[5] (
	.clk(CLK),
	.d(\Mux127~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_5),
	.prn(vcc));
// synopsys translate_off
defparam \pc[5] .is_wysiwyg = "true";
defparam \pc[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y28_N29
dffeas \pc[4] (
	.clk(CLK),
	.d(\Mux128~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_4),
	.prn(vcc));
// synopsys translate_off
defparam \pc[4] .is_wysiwyg = "true";
defparam \pc[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X53_Y29_N25
dffeas \pc[7] (
	.clk(CLK),
	.d(\Mux125~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_7),
	.prn(vcc));
// synopsys translate_off
defparam \pc[7] .is_wysiwyg = "true";
defparam \pc[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N3
dffeas \pc[6] (
	.clk(CLK),
	.d(\Mux126~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_6),
	.prn(vcc));
// synopsys translate_off
defparam \pc[6] .is_wysiwyg = "true";
defparam \pc[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y31_N9
dffeas \pc[9] (
	.clk(CLK),
	.d(\Mux123~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_9),
	.prn(vcc));
// synopsys translate_off
defparam \pc[9] .is_wysiwyg = "true";
defparam \pc[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N25
dffeas \pc[8] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Mux124~1_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_8),
	.prn(vcc));
// synopsys translate_off
defparam \pc[8] .is_wysiwyg = "true";
defparam \pc[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y25_N9
dffeas \pc[11] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Mux121~1_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_11),
	.prn(vcc));
// synopsys translate_off
defparam \pc[11] .is_wysiwyg = "true";
defparam \pc[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y28_N15
dffeas \pc[10] (
	.clk(CLK),
	.d(\Mux122~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_10),
	.prn(vcc));
// synopsys translate_off
defparam \pc[10] .is_wysiwyg = "true";
defparam \pc[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y28_N1
dffeas \pc[13] (
	.clk(CLK),
	.d(\Mux119~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_13),
	.prn(vcc));
// synopsys translate_off
defparam \pc[13] .is_wysiwyg = "true";
defparam \pc[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N13
dffeas \pc[12] (
	.clk(CLK),
	.d(gnd),
	.asdata(\Mux120~1_combout ),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_12),
	.prn(vcc));
// synopsys translate_off
defparam \pc[12] .is_wysiwyg = "true";
defparam \pc[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y26_N15
dffeas \pc[15] (
	.clk(CLK),
	.d(\Mux117~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_15),
	.prn(vcc));
// synopsys translate_off
defparam \pc[15] .is_wysiwyg = "true";
defparam \pc[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y26_N5
dffeas \pc[14] (
	.clk(CLK),
	.d(\Mux118~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_14),
	.prn(vcc));
// synopsys translate_off
defparam \pc[14] .is_wysiwyg = "true";
defparam \pc[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y30_N31
dffeas \pc[23] (
	.clk(CLK),
	.d(\Mux109~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_23),
	.prn(vcc));
// synopsys translate_off
defparam \pc[23] .is_wysiwyg = "true";
defparam \pc[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y30_N29
dffeas \pc[22] (
	.clk(CLK),
	.d(\Mux110~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_22),
	.prn(vcc));
// synopsys translate_off
defparam \pc[22] .is_wysiwyg = "true";
defparam \pc[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y33_N19
dffeas \pc[21] (
	.clk(CLK),
	.d(\Mux111~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_21),
	.prn(vcc));
// synopsys translate_off
defparam \pc[21] .is_wysiwyg = "true";
defparam \pc[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y31_N1
dffeas \pc[29] (
	.clk(CLK),
	.d(\Mux103~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_29),
	.prn(vcc));
// synopsys translate_off
defparam \pc[29] .is_wysiwyg = "true";
defparam \pc[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N29
dffeas \pc[28] (
	.clk(CLK),
	.d(\Mux104~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_28),
	.prn(vcc));
// synopsys translate_off
defparam \pc[28] .is_wysiwyg = "true";
defparam \pc[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N7
dffeas \pc[31] (
	.clk(CLK),
	.d(\Mux101~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_31),
	.prn(vcc));
// synopsys translate_off
defparam \pc[31] .is_wysiwyg = "true";
defparam \pc[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N21
dffeas \pc[30] (
	.clk(CLK),
	.d(\Mux102~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_30),
	.prn(vcc));
// synopsys translate_off
defparam \pc[30] .is_wysiwyg = "true";
defparam \pc[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N25
dffeas \pc[20] (
	.clk(CLK),
	.d(\Mux112~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_20),
	.prn(vcc));
// synopsys translate_off
defparam \pc[20] .is_wysiwyg = "true";
defparam \pc[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N11
dffeas \pc[17] (
	.clk(CLK),
	.d(\Mux115~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_17),
	.prn(vcc));
// synopsys translate_off
defparam \pc[17] .is_wysiwyg = "true";
defparam \pc[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N17
dffeas \pc[16] (
	.clk(CLK),
	.d(\Mux116~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_16),
	.prn(vcc));
// synopsys translate_off
defparam \pc[16] .is_wysiwyg = "true";
defparam \pc[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N19
dffeas \pc[19] (
	.clk(CLK),
	.d(\Mux113~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_19),
	.prn(vcc));
// synopsys translate_off
defparam \pc[19] .is_wysiwyg = "true";
defparam \pc[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y32_N25
dffeas \pc[18] (
	.clk(CLK),
	.d(\Mux114~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_18),
	.prn(vcc));
// synopsys translate_off
defparam \pc[18] .is_wysiwyg = "true";
defparam \pc[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N5
dffeas \pc[25] (
	.clk(CLK),
	.d(\Mux107~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_25),
	.prn(vcc));
// synopsys translate_off
defparam \pc[25] .is_wysiwyg = "true";
defparam \pc[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N31
dffeas \pc[24] (
	.clk(CLK),
	.d(\Mux108~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_24),
	.prn(vcc));
// synopsys translate_off
defparam \pc[24] .is_wysiwyg = "true";
defparam \pc[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N11
dffeas \pc[27] (
	.clk(CLK),
	.d(\Mux105~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_27),
	.prn(vcc));
// synopsys translate_off
defparam \pc[27] .is_wysiwyg = "true";
defparam \pc[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N21
dffeas \pc[26] (
	.clk(CLK),
	.d(\Mux106~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\HU|pc_en~0_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(pc_26),
	.prn(vcc));
// synopsys translate_off
defparam \pc[26] .is_wysiwyg = "true";
defparam \pc[26] .power_up = "low";
// synopsys translate_on

// Location: DDIOOUTCELL_X38_Y0_N4
dffeas \dpif.halt (
	.clk(!CLK),
	.d(\dpif.halt~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(dpifhalt),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt .is_wysiwyg = "true";
defparam \dpif.halt .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N16
cycloneive_lcell_comb \prif.rdat1_mem[21]~0 (
// Equation(s):
// \prif.rdat1_mem[21]~0_combout  = (always1) # ((always1 & ((prifdmemren) # (prifdmemwen))))

	.dataa(prifdmemren),
	.datab(always1),
	.datac(prifdmemwen),
	.datad(\HU|always1~5_combout ),
	.cin(gnd),
	.combout(\prif.rdat1_mem[21]~0_combout ),
	.cout());
// synopsys translate_off
defparam \prif.rdat1_mem[21]~0 .lut_mask = 16'hFFC8;
defparam \prif.rdat1_mem[21]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N13
dffeas \prif.rdat1_mem[1] (
	.clk(CLK),
	.d(\PR|rdat1_mem~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[1] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N31
dffeas \prif.PCScr_mem[0] (
	.clk(CLK),
	.d(\PR|PCScr_mem~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.PCScr_mem [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.PCScr_mem[0] .is_wysiwyg = "true";
defparam \prif.PCScr_mem[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N16
cycloneive_lcell_comb \Mux131~0 (
// Equation(s):
// \Mux131~0_combout  = (\prif.rdat1_mem [1] & !\prif.PCScr_mem [0])

	.dataa(\prif.rdat1_mem [1]),
	.datab(\prif.PCScr_mem [0]),
	.datac(gnd),
	.datad(gnd),
	.cin(gnd),
	.combout(\Mux131~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux131~0 .lut_mask = 16'h2222;
defparam \Mux131~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y26_N5
dffeas \prif.pc_bran_mem[1] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[1] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N19
dffeas \prif.PCScr_mem[1] (
	.clk(CLK),
	.d(\PR|PCScr_mem~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.PCScr_mem [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.PCScr_mem[1] .is_wysiwyg = "true";
defparam \prif.PCScr_mem[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y25_N3
dffeas \prif.zero_flag_mem (
	.clk(CLK),
	.d(\PR|zero_flag_mem~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.zero_flag_mem~q ),
	.prn(vcc));
// synopsys translate_off
defparam \prif.zero_flag_mem .is_wysiwyg = "true";
defparam \prif.zero_flag_mem .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N0
cycloneive_lcell_comb \pc[0]~0 (
// Equation(s):
// \pc[0]~0_combout  = (!\prif.PCScr_mem [1] & ((\Equal1~1_combout  $ (\prif.zero_flag_mem~q )) # (!\prif.PCScr_mem [0])))

	.dataa(\Equal1~1_combout ),
	.datab(\prif.PCScr_mem [1]),
	.datac(\prif.zero_flag_mem~q ),
	.datad(\prif.PCScr_mem [0]),
	.cin(gnd),
	.combout(\pc[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \pc[0]~0 .lut_mask = 16'h1233;
defparam \pc[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N2
cycloneive_lcell_comb \pc[1]~1 (
// Equation(s):
// \pc[1]~1_combout  = (ifid_en & (exmem_en & !\pc[0]~0_combout ))

	.dataa(gnd),
	.datab(\HU|ifid_en~0_combout ),
	.datac(\HU|exmem_en~0_combout ),
	.datad(\pc[0]~0_combout ),
	.cin(gnd),
	.combout(\pc[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \pc[1]~1 .lut_mask = 16'h00C0;
defparam \pc[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N25
dffeas \prif.rdat1_mem[0] (
	.clk(CLK),
	.d(\PR|rdat1_mem~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[0] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N30
cycloneive_lcell_comb \Mux132~0 (
// Equation(s):
// \Mux132~0_combout  = (!\prif.PCScr_mem [0] & \prif.rdat1_mem [0])

	.dataa(gnd),
	.datab(\prif.PCScr_mem [0]),
	.datac(gnd),
	.datad(\prif.rdat1_mem [0]),
	.cin(gnd),
	.combout(\Mux132~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux132~0 .lut_mask = 16'h3300;
defparam \Mux132~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N27
dffeas \prif.pc_bran_mem[0] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[0] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N8
cycloneive_lcell_comb \pc[23]~2 (
// Equation(s):
// \pc[23]~2_combout  = (\prif.PCScr_mem [1] & (((\prif.PCScr_mem [0])))) # (!\prif.PCScr_mem [1] & ((\Equal1~1_combout  $ (\prif.zero_flag_mem~q )) # (!\prif.PCScr_mem [0])))

	.dataa(\Equal1~1_combout ),
	.datab(\prif.PCScr_mem [1]),
	.datac(\prif.zero_flag_mem~q ),
	.datad(\prif.PCScr_mem [0]),
	.cin(gnd),
	.combout(\pc[23]~2_combout ),
	.cout());
// synopsys translate_off
defparam \pc[23]~2 .lut_mask = 16'hDE33;
defparam \pc[23]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N2
cycloneive_lcell_comb \Add3~0 (
// Equation(s):
// \Add3~0_combout  = pc_2 $ (VCC)
// \Add3~1  = CARRY(pc_2)

	.dataa(pc_2),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add3~0_combout ),
	.cout(\Add3~1 ));
// synopsys translate_off
defparam \Add3~0 .lut_mask = 16'h55AA;
defparam \Add3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N4
cycloneive_lcell_comb \Add3~2 (
// Equation(s):
// \Add3~2_combout  = (pc_3 & (!\Add3~1 )) # (!pc_3 & ((\Add3~1 ) # (GND)))
// \Add3~3  = CARRY((!\Add3~1 ) # (!pc_3))

	.dataa(pc_3),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~1 ),
	.combout(\Add3~2_combout ),
	.cout(\Add3~3 ));
// synopsys translate_off
defparam \Add3~2 .lut_mask = 16'h5A5F;
defparam \Add3~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N18
cycloneive_lcell_comb \Mux129~0 (
// Equation(s):
// \Mux129~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & ((\Add3~2_combout ))) # (!\pc[23]~2_combout  & (\prif.pc_bran_mem [3]))))

	.dataa(\prif.pc_bran_mem [3]),
	.datab(\prif.PCScr_mem [1]),
	.datac(\pc[23]~2_combout ),
	.datad(\Add3~2_combout ),
	.cin(gnd),
	.combout(\Mux129~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux129~0 .lut_mask = 16'hF2C2;
defparam \Mux129~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N11
dffeas \prif.instr_mem[1] (
	.clk(CLK),
	.d(\PR|instr_mem~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [1]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[1] .is_wysiwyg = "true";
defparam \prif.instr_mem[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y30_N13
dffeas \prif.rdat1_mem[3] (
	.clk(CLK),
	.d(\PR|rdat1_mem~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[3] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N0
cycloneive_lcell_comb \Mux129~1 (
// Equation(s):
// \Mux129~1_combout  = (\prif.PCScr_mem [1] & ((\Mux129~0_combout  & (\prif.instr_mem [1])) # (!\Mux129~0_combout  & ((\prif.rdat1_mem [3]))))) # (!\prif.PCScr_mem [1] & (\Mux129~0_combout ))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\Mux129~0_combout ),
	.datac(\prif.instr_mem [1]),
	.datad(\prif.rdat1_mem [3]),
	.cin(gnd),
	.combout(\Mux129~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux129~1 .lut_mask = 16'hE6C4;
defparam \Mux129~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N21
dffeas \prif.pc_bran_mem[2] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[2] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N15
dffeas \prif.rdat1_mem[2] (
	.clk(CLK),
	.d(\PR|rdat1_mem~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[2] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N6
cycloneive_lcell_comb \Mux130~0 (
// Equation(s):
// \Mux130~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout ) # (\prif.rdat1_mem [2])))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [2] & (!\pc[23]~2_combout )))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.pc_bran_mem [2]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.rdat1_mem [2]),
	.cin(gnd),
	.combout(\Mux130~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux130~0 .lut_mask = 16'hAEA4;
defparam \Mux130~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N29
dffeas \prif.instr_mem[0] (
	.clk(CLK),
	.d(\PR|instr_mem~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [0]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[0] .is_wysiwyg = "true";
defparam \prif.instr_mem[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N8
cycloneive_lcell_comb \Mux130~1 (
// Equation(s):
// \Mux130~1_combout  = (\Mux130~0_combout  & (((\prif.instr_mem [0])) # (!\pc[23]~2_combout ))) # (!\Mux130~0_combout  & (\pc[23]~2_combout  & ((\Add3~0_combout ))))

	.dataa(\Mux130~0_combout ),
	.datab(\pc[23]~2_combout ),
	.datac(\prif.instr_mem [0]),
	.datad(\Add3~0_combout ),
	.cin(gnd),
	.combout(\Mux130~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux130~1 .lut_mask = 16'hE6A2;
defparam \Mux130~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N21
dffeas \prif.instr_mem[3] (
	.clk(CLK),
	.d(\PR|instr_mem~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [3]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[3] .is_wysiwyg = "true";
defparam \prif.instr_mem[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y28_N21
dffeas \prif.rdat1_mem[5] (
	.clk(CLK),
	.d(\PR|rdat1_mem~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[5] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N6
cycloneive_lcell_comb \Add3~4 (
// Equation(s):
// \Add3~4_combout  = (pc_4 & (\Add3~3  $ (GND))) # (!pc_4 & (!\Add3~3  & VCC))
// \Add3~5  = CARRY((pc_4 & !\Add3~3 ))

	.dataa(pc_4),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~3 ),
	.combout(\Add3~4_combout ),
	.cout(\Add3~5 ));
// synopsys translate_off
defparam \Add3~4 .lut_mask = 16'hA50A;
defparam \Add3~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N8
cycloneive_lcell_comb \Add3~6 (
// Equation(s):
// \Add3~6_combout  = (pc_5 & (!\Add3~5 )) # (!pc_5 & ((\Add3~5 ) # (GND)))
// \Add3~7  = CARRY((!\Add3~5 ) # (!pc_5))

	.dataa(gnd),
	.datab(pc_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~5 ),
	.combout(\Add3~6_combout ),
	.cout(\Add3~7 ));
// synopsys translate_off
defparam \Add3~6 .lut_mask = 16'h3C3F;
defparam \Add3~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X54_Y31_N23
dffeas \prif.pc_bran_mem[5] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~4_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[5] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N0
cycloneive_lcell_comb \Mux127~0 (
// Equation(s):
// \Mux127~0_combout  = (\prif.PCScr_mem [1] & (\pc[23]~2_combout )) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & (\Add3~6_combout )) # (!\pc[23]~2_combout  & ((\prif.pc_bran_mem [5])))))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\pc[23]~2_combout ),
	.datac(\Add3~6_combout ),
	.datad(\prif.pc_bran_mem [5]),
	.cin(gnd),
	.combout(\Mux127~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux127~0 .lut_mask = 16'hD9C8;
defparam \Mux127~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N22
cycloneive_lcell_comb \Mux127~1 (
// Equation(s):
// \Mux127~1_combout  = (\prif.PCScr_mem [1] & ((\Mux127~0_combout  & (\prif.instr_mem [3])) # (!\Mux127~0_combout  & ((\prif.rdat1_mem [5]))))) # (!\prif.PCScr_mem [1] & (((\Mux127~0_combout ))))

	.dataa(\prif.instr_mem [3]),
	.datab(\prif.rdat1_mem [5]),
	.datac(\prif.PCScr_mem [1]),
	.datad(\Mux127~0_combout ),
	.cin(gnd),
	.combout(\Mux127~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux127~1 .lut_mask = 16'hAFC0;
defparam \Mux127~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y30_N17
dffeas \prif.instr_mem[2] (
	.clk(CLK),
	.d(\PR|instr_mem~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [2]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[2] .is_wysiwyg = "true";
defparam \prif.instr_mem[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N9
dffeas \prif.rdat1_mem[4] (
	.clk(CLK),
	.d(\PR|rdat1_mem~5_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[4] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N24
cycloneive_lcell_comb \Mux128~0 (
// Equation(s):
// \Mux128~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout ) # (\prif.rdat1_mem [4])))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [4] & (!\pc[23]~2_combout )))

	.dataa(\prif.pc_bran_mem [4]),
	.datab(\prif.PCScr_mem [1]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.rdat1_mem [4]),
	.cin(gnd),
	.combout(\Mux128~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux128~0 .lut_mask = 16'hCEC2;
defparam \Mux128~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N28
cycloneive_lcell_comb \Mux128~1 (
// Equation(s):
// \Mux128~1_combout  = (\Mux128~0_combout  & ((\prif.instr_mem [2]) # ((!\pc[23]~2_combout )))) # (!\Mux128~0_combout  & (((\Add3~4_combout  & \pc[23]~2_combout ))))

	.dataa(\prif.instr_mem [2]),
	.datab(\Mux128~0_combout ),
	.datac(\Add3~4_combout ),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux128~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux128~1 .lut_mask = 16'hB8CC;
defparam \Mux128~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N19
dffeas \prif.rdat1_mem[7] (
	.clk(CLK),
	.d(\PR|rdat1_mem~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[7] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N31
dffeas \prif.pc_bran_mem[7] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[7] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N10
cycloneive_lcell_comb \Add3~8 (
// Equation(s):
// \Add3~8_combout  = (pc_6 & (\Add3~7  $ (GND))) # (!pc_6 & (!\Add3~7  & VCC))
// \Add3~9  = CARRY((pc_6 & !\Add3~7 ))

	.dataa(gnd),
	.datab(pc_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~7 ),
	.combout(\Add3~8_combout ),
	.cout(\Add3~9 ));
// synopsys translate_off
defparam \Add3~8 .lut_mask = 16'hC30C;
defparam \Add3~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N12
cycloneive_lcell_comb \Add3~10 (
// Equation(s):
// \Add3~10_combout  = (pc_7 & (!\Add3~9 )) # (!pc_7 & ((\Add3~9 ) # (GND)))
// \Add3~11  = CARRY((!\Add3~9 ) # (!pc_7))

	.dataa(pc_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~9 ),
	.combout(\Add3~10_combout ),
	.cout(\Add3~11 ));
// synopsys translate_off
defparam \Add3~10 .lut_mask = 16'h5A5F;
defparam \Add3~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N26
cycloneive_lcell_comb \Mux125~0 (
// Equation(s):
// \Mux125~0_combout  = (\pc[23]~2_combout  & ((\prif.PCScr_mem [1]) # ((\Add3~10_combout )))) # (!\pc[23]~2_combout  & (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [7])))

	.dataa(\pc[23]~2_combout ),
	.datab(\prif.PCScr_mem [1]),
	.datac(\prif.pc_bran_mem [7]),
	.datad(\Add3~10_combout ),
	.cin(gnd),
	.combout(\Mux125~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux125~0 .lut_mask = 16'hBA98;
defparam \Mux125~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N7
dffeas \prif.instr_mem[5] (
	.clk(CLK),
	.d(\PR|instr_mem~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [5]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[5] .is_wysiwyg = "true";
defparam \prif.instr_mem[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N24
cycloneive_lcell_comb \Mux125~1 (
// Equation(s):
// \Mux125~1_combout  = (\Mux125~0_combout  & (((\prif.instr_mem [5]) # (!\prif.PCScr_mem [1])))) # (!\Mux125~0_combout  & (\prif.rdat1_mem [7] & ((\prif.PCScr_mem [1]))))

	.dataa(\prif.rdat1_mem [7]),
	.datab(\Mux125~0_combout ),
	.datac(\prif.instr_mem [5]),
	.datad(\prif.PCScr_mem [1]),
	.cin(gnd),
	.combout(\Mux125~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux125~1 .lut_mask = 16'hE2CC;
defparam \Mux125~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N13
dffeas \prif.instr_mem[4] (
	.clk(CLK),
	.d(\PR|instr_mem~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [4]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[4] .is_wysiwyg = "true";
defparam \prif.instr_mem[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N7
dffeas \prif.pc_bran_mem[6] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[6] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N29
dffeas \prif.rdat1_mem[6] (
	.clk(CLK),
	.d(\PR|rdat1_mem~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[6] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N18
cycloneive_lcell_comb \Mux126~0 (
// Equation(s):
// \Mux126~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout ) # (\prif.rdat1_mem [6])))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [6] & (!\pc[23]~2_combout )))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.pc_bran_mem [6]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.rdat1_mem [6]),
	.cin(gnd),
	.combout(\Mux126~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux126~0 .lut_mask = 16'hAEA4;
defparam \Mux126~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N2
cycloneive_lcell_comb \Mux126~1 (
// Equation(s):
// \Mux126~1_combout  = (\Mux126~0_combout  & ((\prif.instr_mem [4]) # ((!\pc[23]~2_combout )))) # (!\Mux126~0_combout  & (((\pc[23]~2_combout  & \Add3~8_combout ))))

	.dataa(\prif.instr_mem [4]),
	.datab(\Mux126~0_combout ),
	.datac(\pc[23]~2_combout ),
	.datad(\Add3~8_combout ),
	.cin(gnd),
	.combout(\Mux126~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux126~1 .lut_mask = 16'hBC8C;
defparam \Mux126~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y31_N11
dffeas \prif.instr_mem[7] (
	.clk(CLK),
	.d(\PR|instr_mem~6_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [7]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[7] .is_wysiwyg = "true";
defparam \prif.instr_mem[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y31_N17
dffeas \prif.rdat1_mem[9] (
	.clk(CLK),
	.d(\PR|rdat1_mem~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[9] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N13
dffeas \prif.pc_bran_mem[9] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[9] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N10
cycloneive_lcell_comb \Mux123~0 (
// Equation(s):
// \Mux123~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & (\Add3~14_combout )) # (!\pc[23]~2_combout  & ((\prif.pc_bran_mem [9])))))

	.dataa(\Add3~14_combout ),
	.datab(\prif.PCScr_mem [1]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.pc_bran_mem [9]),
	.cin(gnd),
	.combout(\Mux123~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux123~0 .lut_mask = 16'hE3E0;
defparam \Mux123~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N8
cycloneive_lcell_comb \Mux123~1 (
// Equation(s):
// \Mux123~1_combout  = (\prif.PCScr_mem [1] & ((\Mux123~0_combout  & (\prif.instr_mem [7])) # (!\Mux123~0_combout  & ((\prif.rdat1_mem [9]))))) # (!\prif.PCScr_mem [1] & (((\Mux123~0_combout ))))

	.dataa(\prif.instr_mem [7]),
	.datab(\prif.rdat1_mem [9]),
	.datac(\prif.PCScr_mem [1]),
	.datad(\Mux123~0_combout ),
	.cin(gnd),
	.combout(\Mux123~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux123~1 .lut_mask = 16'hAFC0;
defparam \Mux123~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N14
cycloneive_lcell_comb \Add3~12 (
// Equation(s):
// \Add3~12_combout  = (pc_8 & (\Add3~11  $ (GND))) # (!pc_8 & (!\Add3~11  & VCC))
// \Add3~13  = CARRY((pc_8 & !\Add3~11 ))

	.dataa(gnd),
	.datab(pc_8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~11 ),
	.combout(\Add3~12_combout ),
	.cout(\Add3~13 ));
// synopsys translate_off
defparam \Add3~12 .lut_mask = 16'hC30C;
defparam \Add3~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X57_Y32_N19
dffeas \prif.instr_mem[6] (
	.clk(CLK),
	.d(\PR|instr_mem~7_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [6]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[6] .is_wysiwyg = "true";
defparam \prif.instr_mem[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N17
dffeas \prif.pc_bran_mem[8] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[8] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N0
cycloneive_lcell_comb \Mux124~0 (
// Equation(s):
// \Mux124~0_combout  = (\prif.PCScr_mem [1] & ((\prif.rdat1_mem [8]) # ((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & (((!\pc[23]~2_combout  & \prif.pc_bran_mem [8]))))

	.dataa(\prif.rdat1_mem [8]),
	.datab(\prif.PCScr_mem [1]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.pc_bran_mem [8]),
	.cin(gnd),
	.combout(\Mux124~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux124~0 .lut_mask = 16'hCBC8;
defparam \Mux124~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N0
cycloneive_lcell_comb \Mux124~1 (
// Equation(s):
// \Mux124~1_combout  = (\pc[23]~2_combout  & ((\Mux124~0_combout  & ((\prif.instr_mem [6]))) # (!\Mux124~0_combout  & (\Add3~12_combout )))) # (!\pc[23]~2_combout  & (((\Mux124~0_combout ))))

	.dataa(\pc[23]~2_combout ),
	.datab(\Add3~12_combout ),
	.datac(\prif.instr_mem [6]),
	.datad(\Mux124~0_combout ),
	.cin(gnd),
	.combout(\Mux124~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux124~1 .lut_mask = 16'hF588;
defparam \Mux124~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y28_N13
dffeas \prif.instr_mem[9] (
	.clk(CLK),
	.d(\PR|instr_mem~8_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [9]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[9] .is_wysiwyg = "true";
defparam \prif.instr_mem[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N25
dffeas \prif.pc_bran_mem[11] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[11] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N18
cycloneive_lcell_comb \Add3~16 (
// Equation(s):
// \Add3~16_combout  = (pc_10 & (\Add3~15  $ (GND))) # (!pc_10 & (!\Add3~15  & VCC))
// \Add3~17  = CARRY((pc_10 & !\Add3~15 ))

	.dataa(gnd),
	.datab(pc_10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~15 ),
	.combout(\Add3~16_combout ),
	.cout(\Add3~17 ));
// synopsys translate_off
defparam \Add3~16 .lut_mask = 16'hC30C;
defparam \Add3~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N20
cycloneive_lcell_comb \Add3~18 (
// Equation(s):
// \Add3~18_combout  = (pc_11 & (!\Add3~17 )) # (!pc_11 & ((\Add3~17 ) # (GND)))
// \Add3~19  = CARRY((!\Add3~17 ) # (!pc_11))

	.dataa(gnd),
	.datab(pc_11),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~17 ),
	.combout(\Add3~18_combout ),
	.cout(\Add3~19 ));
// synopsys translate_off
defparam \Add3~18 .lut_mask = 16'h3C3F;
defparam \Add3~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N22
cycloneive_lcell_comb \Mux121~0 (
// Equation(s):
// \Mux121~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & ((\Add3~18_combout ))) # (!\pc[23]~2_combout  & (\prif.pc_bran_mem [11]))))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.pc_bran_mem [11]),
	.datac(\Add3~18_combout ),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux121~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux121~0 .lut_mask = 16'hFA44;
defparam \Mux121~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y28_N3
dffeas \prif.rdat1_mem[11] (
	.clk(CLK),
	.d(\PR|rdat1_mem~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[11] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N10
cycloneive_lcell_comb \Mux121~1 (
// Equation(s):
// \Mux121~1_combout  = (\Mux121~0_combout  & ((\prif.instr_mem [9]) # ((!\prif.PCScr_mem [1])))) # (!\Mux121~0_combout  & (((\prif.PCScr_mem [1] & \prif.rdat1_mem [11]))))

	.dataa(\prif.instr_mem [9]),
	.datab(\Mux121~0_combout ),
	.datac(\prif.PCScr_mem [1]),
	.datad(\prif.rdat1_mem [11]),
	.cin(gnd),
	.combout(\Mux121~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux121~1 .lut_mask = 16'hBC8C;
defparam \Mux121~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y28_N7
dffeas \prif.instr_mem[8] (
	.clk(CLK),
	.d(\PR|instr_mem~9_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [8]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[8] .is_wysiwyg = "true";
defparam \prif.instr_mem[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y28_N17
dffeas \prif.pc_bran_mem[10] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[10] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N4
cycloneive_lcell_comb \Mux122~0 (
// Equation(s):
// \Mux122~0_combout  = (\prif.PCScr_mem [1] & ((\prif.rdat1_mem [10]) # ((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & (((\prif.pc_bran_mem [10] & !\pc[23]~2_combout ))))

	.dataa(\prif.rdat1_mem [10]),
	.datab(\prif.pc_bran_mem [10]),
	.datac(\prif.PCScr_mem [1]),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux122~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux122~0 .lut_mask = 16'hF0AC;
defparam \Mux122~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N14
cycloneive_lcell_comb \Mux122~1 (
// Equation(s):
// \Mux122~1_combout  = (\Mux122~0_combout  & ((\prif.instr_mem [8]) # ((!\pc[23]~2_combout )))) # (!\Mux122~0_combout  & (((\Add3~16_combout  & \pc[23]~2_combout ))))

	.dataa(\prif.instr_mem [8]),
	.datab(\Mux122~0_combout ),
	.datac(\Add3~16_combout ),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux122~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux122~1 .lut_mask = 16'hB8CC;
defparam \Mux122~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N22
cycloneive_lcell_comb \Add3~20 (
// Equation(s):
// \Add3~20_combout  = (pc_12 & (\Add3~19  $ (GND))) # (!pc_12 & (!\Add3~19  & VCC))
// \Add3~21  = CARRY((pc_12 & !\Add3~19 ))

	.dataa(gnd),
	.datab(pc_12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~19 ),
	.combout(\Add3~20_combout ),
	.cout(\Add3~21 ));
// synopsys translate_off
defparam \Add3~20 .lut_mask = 16'hC30C;
defparam \Add3~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N24
cycloneive_lcell_comb \Add3~22 (
// Equation(s):
// \Add3~22_combout  = (pc_13 & (!\Add3~21 )) # (!pc_13 & ((\Add3~21 ) # (GND)))
// \Add3~23  = CARRY((!\Add3~21 ) # (!pc_13))

	.dataa(gnd),
	.datab(pc_13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~21 ),
	.combout(\Add3~22_combout ),
	.cout(\Add3~23 ));
// synopsys translate_off
defparam \Add3~22 .lut_mask = 16'h3C3F;
defparam \Add3~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X58_Y28_N25
dffeas \prif.pc_bran_mem[13] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[13] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N26
cycloneive_lcell_comb \Mux119~0 (
// Equation(s):
// \Mux119~0_combout  = (\pc[23]~2_combout  & ((\Add3~22_combout ) # ((\prif.PCScr_mem [1])))) # (!\pc[23]~2_combout  & (((!\prif.PCScr_mem [1] & \prif.pc_bran_mem [13]))))

	.dataa(\pc[23]~2_combout ),
	.datab(\Add3~22_combout ),
	.datac(\prif.PCScr_mem [1]),
	.datad(\prif.pc_bran_mem [13]),
	.cin(gnd),
	.combout(\Mux119~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux119~0 .lut_mask = 16'hADA8;
defparam \Mux119~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y28_N31
dffeas \prif.instr_mem[11] (
	.clk(CLK),
	.d(\PR|instr_mem~10_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [11]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[11] .is_wysiwyg = "true";
defparam \prif.instr_mem[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N11
dffeas \prif.rdat1_mem[13] (
	.clk(CLK),
	.d(\PR|rdat1_mem~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[13] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N0
cycloneive_lcell_comb \Mux119~1 (
// Equation(s):
// \Mux119~1_combout  = (\Mux119~0_combout  & (((\prif.instr_mem [11])) # (!\prif.PCScr_mem [1]))) # (!\Mux119~0_combout  & (\prif.PCScr_mem [1] & ((\prif.rdat1_mem [13]))))

	.dataa(\Mux119~0_combout ),
	.datab(\prif.PCScr_mem [1]),
	.datac(\prif.instr_mem [11]),
	.datad(\prif.rdat1_mem [13]),
	.cin(gnd),
	.combout(\Mux119~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux119~1 .lut_mask = 16'hE6A2;
defparam \Mux119~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N1
dffeas \prif.instr_mem[10] (
	.clk(CLK),
	.d(\PR|instr_mem~11_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [10]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[10] .is_wysiwyg = "true";
defparam \prif.instr_mem[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N15
dffeas \prif.pc_bran_mem[12] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[12] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N25
dffeas \prif.rdat1_mem[12] (
	.clk(CLK),
	.d(\PR|rdat1_mem~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[12] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N18
cycloneive_lcell_comb \Mux120~0 (
// Equation(s):
// \Mux120~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout ) # (\prif.rdat1_mem [12])))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [12] & (!\pc[23]~2_combout )))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.pc_bran_mem [12]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.rdat1_mem [12]),
	.cin(gnd),
	.combout(\Mux120~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux120~0 .lut_mask = 16'hAEA4;
defparam \Mux120~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N4
cycloneive_lcell_comb \Mux120~1 (
// Equation(s):
// \Mux120~1_combout  = (\pc[23]~2_combout  & ((\Mux120~0_combout  & (\prif.instr_mem [10])) # (!\Mux120~0_combout  & ((\Add3~20_combout ))))) # (!\pc[23]~2_combout  & (((\Mux120~0_combout ))))

	.dataa(\pc[23]~2_combout ),
	.datab(\prif.instr_mem [10]),
	.datac(\Add3~20_combout ),
	.datad(\Mux120~0_combout ),
	.cin(gnd),
	.combout(\Mux120~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux120~1 .lut_mask = 16'hDDA0;
defparam \Mux120~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y26_N23
dffeas \prif.rdat1_mem[15] (
	.clk(CLK),
	.d(\PR|rdat1_mem~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[15] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y26_N1
dffeas \prif.instr_mem[13] (
	.clk(CLK),
	.d(\PR|instr_mem~12_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [13]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[13] .is_wysiwyg = "true";
defparam \prif.instr_mem[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N7
dffeas \prif.pc_bran_mem[15] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[15] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N26
cycloneive_lcell_comb \Add3~24 (
// Equation(s):
// \Add3~24_combout  = (pc_14 & (\Add3~23  $ (GND))) # (!pc_14 & (!\Add3~23  & VCC))
// \Add3~25  = CARRY((pc_14 & !\Add3~23 ))

	.dataa(pc_14),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~23 ),
	.combout(\Add3~24_combout ),
	.cout(\Add3~25 ));
// synopsys translate_off
defparam \Add3~24 .lut_mask = 16'hA50A;
defparam \Add3~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N28
cycloneive_lcell_comb \Add3~26 (
// Equation(s):
// \Add3~26_combout  = (pc_15 & (!\Add3~25 )) # (!pc_15 & ((\Add3~25 ) # (GND)))
// \Add3~27  = CARRY((!\Add3~25 ) # (!pc_15))

	.dataa(pc_15),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~25 ),
	.combout(\Add3~26_combout ),
	.cout(\Add3~27 ));
// synopsys translate_off
defparam \Add3~26 .lut_mask = 16'h5A5F;
defparam \Add3~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N26
cycloneive_lcell_comb \Mux117~0 (
// Equation(s):
// \Mux117~0_combout  = (\prif.PCScr_mem [1] & (\pc[23]~2_combout )) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & ((\Add3~26_combout ))) # (!\pc[23]~2_combout  & (\prif.pc_bran_mem [15]))))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\pc[23]~2_combout ),
	.datac(\prif.pc_bran_mem [15]),
	.datad(\Add3~26_combout ),
	.cin(gnd),
	.combout(\Mux117~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux117~0 .lut_mask = 16'hDC98;
defparam \Mux117~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N14
cycloneive_lcell_comb \Mux117~1 (
// Equation(s):
// \Mux117~1_combout  = (\Mux117~0_combout  & (((\prif.instr_mem [13]) # (!\prif.PCScr_mem [1])))) # (!\Mux117~0_combout  & (\prif.rdat1_mem [15] & ((\prif.PCScr_mem [1]))))

	.dataa(\prif.rdat1_mem [15]),
	.datab(\prif.instr_mem [13]),
	.datac(\Mux117~0_combout ),
	.datad(\prif.PCScr_mem [1]),
	.cin(gnd),
	.combout(\Mux117~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux117~1 .lut_mask = 16'hCAF0;
defparam \Mux117~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N3
dffeas \prif.instr_mem[12] (
	.clk(CLK),
	.d(\PR|instr_mem~13_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [12]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[12] .is_wysiwyg = "true";
defparam \prif.instr_mem[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N21
dffeas \prif.pc_bran_mem[14] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[14] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N7
dffeas \prif.rdat1_mem[14] (
	.clk(CLK),
	.d(\PR|rdat1_mem~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[14] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N22
cycloneive_lcell_comb \Mux118~0 (
// Equation(s):
// \Mux118~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout ) # (\prif.rdat1_mem [14])))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [14] & (!\pc[23]~2_combout )))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.pc_bran_mem [14]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.rdat1_mem [14]),
	.cin(gnd),
	.combout(\Mux118~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux118~0 .lut_mask = 16'hAEA4;
defparam \Mux118~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N4
cycloneive_lcell_comb \Mux118~1 (
// Equation(s):
// \Mux118~1_combout  = (\pc[23]~2_combout  & ((\Mux118~0_combout  & ((\prif.instr_mem [12]))) # (!\Mux118~0_combout  & (\Add3~24_combout )))) # (!\pc[23]~2_combout  & (((\Mux118~0_combout ))))

	.dataa(\Add3~24_combout ),
	.datab(\prif.instr_mem [12]),
	.datac(\pc[23]~2_combout ),
	.datad(\Mux118~0_combout ),
	.cin(gnd),
	.combout(\Mux118~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux118~1 .lut_mask = 16'hCFA0;
defparam \Mux118~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N9
dffeas \prif.rdat1_mem[23] (
	.clk(CLK),
	.d(\PR|rdat1_mem~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[23] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y30_N17
dffeas \prif.instr_mem[21] (
	.clk(CLK),
	.d(\PR|instr_mem~14_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[21] .is_wysiwyg = "true";
defparam \prif.instr_mem[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N30
cycloneive_lcell_comb \Add3~28 (
// Equation(s):
// \Add3~28_combout  = (pc_16 & (\Add3~27  $ (GND))) # (!pc_16 & (!\Add3~27  & VCC))
// \Add3~29  = CARRY((pc_16 & !\Add3~27 ))

	.dataa(gnd),
	.datab(pc_16),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~27 ),
	.combout(\Add3~28_combout ),
	.cout(\Add3~29 ));
// synopsys translate_off
defparam \Add3~28 .lut_mask = 16'hC30C;
defparam \Add3~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N2
cycloneive_lcell_comb \Add3~32 (
// Equation(s):
// \Add3~32_combout  = (pc_18 & (\Add3~31  $ (GND))) # (!pc_18 & (!\Add3~31  & VCC))
// \Add3~33  = CARRY((pc_18 & !\Add3~31 ))

	.dataa(gnd),
	.datab(pc_18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~31 ),
	.combout(\Add3~32_combout ),
	.cout(\Add3~33 ));
// synopsys translate_off
defparam \Add3~32 .lut_mask = 16'hC30C;
defparam \Add3~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N6
cycloneive_lcell_comb \Add3~36 (
// Equation(s):
// \Add3~36_combout  = (pc_20 & (\Add3~35  $ (GND))) # (!pc_20 & (!\Add3~35  & VCC))
// \Add3~37  = CARRY((pc_20 & !\Add3~35 ))

	.dataa(pc_20),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~35 ),
	.combout(\Add3~36_combout ),
	.cout(\Add3~37 ));
// synopsys translate_off
defparam \Add3~36 .lut_mask = 16'hA50A;
defparam \Add3~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N8
cycloneive_lcell_comb \Add3~38 (
// Equation(s):
// \Add3~38_combout  = (pc_21 & (!\Add3~37 )) # (!pc_21 & ((\Add3~37 ) # (GND)))
// \Add3~39  = CARRY((!\Add3~37 ) # (!pc_21))

	.dataa(gnd),
	.datab(pc_21),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~37 ),
	.combout(\Add3~38_combout ),
	.cout(\Add3~39 ));
// synopsys translate_off
defparam \Add3~38 .lut_mask = 16'h3C3F;
defparam \Add3~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N10
cycloneive_lcell_comb \Add3~40 (
// Equation(s):
// \Add3~40_combout  = (pc_22 & (\Add3~39  $ (GND))) # (!pc_22 & (!\Add3~39  & VCC))
// \Add3~41  = CARRY((pc_22 & !\Add3~39 ))

	.dataa(gnd),
	.datab(pc_22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~39 ),
	.combout(\Add3~40_combout ),
	.cout(\Add3~41 ));
// synopsys translate_off
defparam \Add3~40 .lut_mask = 16'hC30C;
defparam \Add3~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N12
cycloneive_lcell_comb \Add3~42 (
// Equation(s):
// \Add3~42_combout  = (pc_23 & (!\Add3~41 )) # (!pc_23 & ((\Add3~41 ) # (GND)))
// \Add3~43  = CARRY((!\Add3~41 ) # (!pc_23))

	.dataa(pc_23),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~41 ),
	.combout(\Add3~42_combout ),
	.cout(\Add3~43 ));
// synopsys translate_off
defparam \Add3~42 .lut_mask = 16'h5A5F;
defparam \Add3~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N12
cycloneive_lcell_comb \Mux109~0 (
// Equation(s):
// \Mux109~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & ((\Add3~42_combout ))) # (!\pc[23]~2_combout  & (\prif.pc_bran_mem [23]))))

	.dataa(\prif.pc_bran_mem [23]),
	.datab(\Add3~42_combout ),
	.datac(\prif.PCScr_mem [1]),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux109~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux109~0 .lut_mask = 16'hFC0A;
defparam \Mux109~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N30
cycloneive_lcell_comb \Mux109~1 (
// Equation(s):
// \Mux109~1_combout  = (\prif.PCScr_mem [1] & ((\Mux109~0_combout  & ((\prif.instr_mem [21]))) # (!\Mux109~0_combout  & (\prif.rdat1_mem [23])))) # (!\prif.PCScr_mem [1] & (((\Mux109~0_combout ))))

	.dataa(\prif.rdat1_mem [23]),
	.datab(\prif.PCScr_mem [1]),
	.datac(\prif.instr_mem [21]),
	.datad(\Mux109~0_combout ),
	.cin(gnd),
	.combout(\Mux109~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux109~1 .lut_mask = 16'hF388;
defparam \Mux109~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N21
dffeas \prif.rdat1_mem[22] (
	.clk(CLK),
	.d(\PR|rdat1_mem~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[22] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N30
cycloneive_lcell_comb \Mux110~0 (
// Equation(s):
// \Mux110~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout ) # (\prif.rdat1_mem [22])))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [22] & (!\pc[23]~2_combout )))

	.dataa(\prif.pc_bran_mem [22]),
	.datab(\prif.PCScr_mem [1]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.rdat1_mem [22]),
	.cin(gnd),
	.combout(\Mux110~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux110~0 .lut_mask = 16'hCEC2;
defparam \Mux110~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y28_N9
dffeas \prif.instr_mem[20] (
	.clk(CLK),
	.d(\PR|instr_mem~15_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[20] .is_wysiwyg = "true";
defparam \prif.instr_mem[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N28
cycloneive_lcell_comb \Mux110~1 (
// Equation(s):
// \Mux110~1_combout  = (\Mux110~0_combout  & (((\prif.instr_mem [20]) # (!\pc[23]~2_combout )))) # (!\Mux110~0_combout  & (\Add3~40_combout  & ((\pc[23]~2_combout ))))

	.dataa(\Mux110~0_combout ),
	.datab(\Add3~40_combout ),
	.datac(\prif.instr_mem [20]),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux110~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux110~1 .lut_mask = 16'hE4AA;
defparam \Mux110~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y33_N1
dffeas \prif.instr_mem[19] (
	.clk(CLK),
	.d(\PR|instr_mem~16_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[19] .is_wysiwyg = "true";
defparam \prif.instr_mem[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N17
dffeas \prif.rdat1_mem[21] (
	.clk(CLK),
	.d(\PR|rdat1_mem~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[21] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N19
dffeas \prif.pc_bran_mem[21] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [21]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[21] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N24
cycloneive_lcell_comb \Mux111~0 (
// Equation(s):
// \Mux111~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & ((\Add3~38_combout ))) # (!\pc[23]~2_combout  & (\prif.pc_bran_mem [21]))))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.pc_bran_mem [21]),
	.datac(\pc[23]~2_combout ),
	.datad(\Add3~38_combout ),
	.cin(gnd),
	.combout(\Mux111~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux111~0 .lut_mask = 16'hF4A4;
defparam \Mux111~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N18
cycloneive_lcell_comb \Mux111~1 (
// Equation(s):
// \Mux111~1_combout  = (\prif.PCScr_mem [1] & ((\Mux111~0_combout  & (\prif.instr_mem [19])) # (!\Mux111~0_combout  & ((\prif.rdat1_mem [21]))))) # (!\prif.PCScr_mem [1] & (((\Mux111~0_combout ))))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.instr_mem [19]),
	.datac(\prif.rdat1_mem [21]),
	.datad(\Mux111~0_combout ),
	.cin(gnd),
	.combout(\Mux111~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux111~1 .lut_mask = 16'hDDA0;
defparam \Mux111~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N25
dffeas \prif.rdat1_mem[29] (
	.clk(CLK),
	.d(\PR|rdat1_mem~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[29] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N20
cycloneive_lcell_comb \Mux103~0 (
// Equation(s):
// \Mux103~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout ) # (\prif.rdat1_mem [29])))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [29] & (!\pc[23]~2_combout )))

	.dataa(\prif.pc_bran_mem [29]),
	.datab(\prif.PCScr_mem [1]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.rdat1_mem [29]),
	.cin(gnd),
	.combout(\Mux103~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux103~0 .lut_mask = 16'hCEC2;
defparam \Mux103~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y31_N7
dffeas \prif.pc_mem[29] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[29]~0_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [29]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[29] .is_wysiwyg = "true";
defparam \prif.pc_mem[29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N14
cycloneive_lcell_comb \Add3~44 (
// Equation(s):
// \Add3~44_combout  = (pc_24 & (\Add3~43  $ (GND))) # (!pc_24 & (!\Add3~43  & VCC))
// \Add3~45  = CARRY((pc_24 & !\Add3~43 ))

	.dataa(gnd),
	.datab(pc_24),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~43 ),
	.combout(\Add3~44_combout ),
	.cout(\Add3~45 ));
// synopsys translate_off
defparam \Add3~44 .lut_mask = 16'hC30C;
defparam \Add3~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N18
cycloneive_lcell_comb \Add3~48 (
// Equation(s):
// \Add3~48_combout  = (pc_26 & (\Add3~47  $ (GND))) # (!pc_26 & (!\Add3~47  & VCC))
// \Add3~49  = CARRY((pc_26 & !\Add3~47 ))

	.dataa(pc_26),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~47 ),
	.combout(\Add3~48_combout ),
	.cout(\Add3~49 ));
// synopsys translate_off
defparam \Add3~48 .lut_mask = 16'hA50A;
defparam \Add3~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N20
cycloneive_lcell_comb \Add3~50 (
// Equation(s):
// \Add3~50_combout  = (pc_27 & (!\Add3~49 )) # (!pc_27 & ((\Add3~49 ) # (GND)))
// \Add3~51  = CARRY((!\Add3~49 ) # (!pc_27))

	.dataa(gnd),
	.datab(pc_27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~49 ),
	.combout(\Add3~50_combout ),
	.cout(\Add3~51 ));
// synopsys translate_off
defparam \Add3~50 .lut_mask = 16'h3C3F;
defparam \Add3~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N22
cycloneive_lcell_comb \Add3~52 (
// Equation(s):
// \Add3~52_combout  = (pc_28 & (\Add3~51  $ (GND))) # (!pc_28 & (!\Add3~51  & VCC))
// \Add3~53  = CARRY((pc_28 & !\Add3~51 ))

	.dataa(gnd),
	.datab(pc_28),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~51 ),
	.combout(\Add3~52_combout ),
	.cout(\Add3~53 ));
// synopsys translate_off
defparam \Add3~52 .lut_mask = 16'hC30C;
defparam \Add3~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N24
cycloneive_lcell_comb \Add3~54 (
// Equation(s):
// \Add3~54_combout  = (pc_29 & (!\Add3~53 )) # (!pc_29 & ((\Add3~53 ) # (GND)))
// \Add3~55  = CARRY((!\Add3~53 ) # (!pc_29))

	.dataa(gnd),
	.datab(pc_29),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~53 ),
	.combout(\Add3~54_combout ),
	.cout(\Add3~55 ));
// synopsys translate_off
defparam \Add3~54 .lut_mask = 16'h3C3F;
defparam \Add3~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y31_N0
cycloneive_lcell_comb \Mux103~1 (
// Equation(s):
// \Mux103~1_combout  = (\Mux103~0_combout  & ((\prif.pc_mem [29]) # ((!\pc[23]~2_combout )))) # (!\Mux103~0_combout  & (((\Add3~54_combout  & \pc[23]~2_combout ))))

	.dataa(\Mux103~0_combout ),
	.datab(\prif.pc_mem [29]),
	.datac(\Add3~54_combout ),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux103~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux103~1 .lut_mask = 16'hD8AA;
defparam \Mux103~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N5
dffeas \prif.pc_mem[28] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[28]~1_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[28] .is_wysiwyg = "true";
defparam \prif.pc_mem[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N5
dffeas \prif.pc_bran_mem[28] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[28] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N3
dffeas \prif.rdat1_mem[28] (
	.clk(CLK),
	.d(\PR|rdat1_mem~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [28]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[28] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N22
cycloneive_lcell_comb \Mux104~0 (
// Equation(s):
// \Mux104~0_combout  = (\pc[23]~2_combout  & (((\prif.PCScr_mem [1])))) # (!\pc[23]~2_combout  & ((\prif.PCScr_mem [1] & ((\prif.rdat1_mem [28]))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [28]))))

	.dataa(\pc[23]~2_combout ),
	.datab(\prif.pc_bran_mem [28]),
	.datac(\prif.PCScr_mem [1]),
	.datad(\prif.rdat1_mem [28]),
	.cin(gnd),
	.combout(\Mux104~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux104~0 .lut_mask = 16'hF4A4;
defparam \Mux104~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N28
cycloneive_lcell_comb \Mux104~1 (
// Equation(s):
// \Mux104~1_combout  = (\Mux104~0_combout  & (((\prif.pc_mem [28]) # (!\pc[23]~2_combout )))) # (!\Mux104~0_combout  & (\Add3~52_combout  & ((\pc[23]~2_combout ))))

	.dataa(\Add3~52_combout ),
	.datab(\prif.pc_mem [28]),
	.datac(\Mux104~0_combout ),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux104~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux104~1 .lut_mask = 16'hCAF0;
defparam \Mux104~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N26
cycloneive_lcell_comb \Add3~56 (
// Equation(s):
// \Add3~56_combout  = (pc_30 & (\Add3~55  $ (GND))) # (!pc_30 & (!\Add3~55  & VCC))
// \Add3~57  = CARRY((pc_30 & !\Add3~55 ))

	.dataa(gnd),
	.datab(pc_30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add3~55 ),
	.combout(\Add3~56_combout ),
	.cout(\Add3~57 ));
// synopsys translate_off
defparam \Add3~56 .lut_mask = 16'hC30C;
defparam \Add3~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y30_N28
cycloneive_lcell_comb \Add3~58 (
// Equation(s):
// \Add3~58_combout  = pc_31 $ (\Add3~57 )

	.dataa(gnd),
	.datab(pc_31),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add3~57 ),
	.combout(\Add3~58_combout ),
	.cout());
// synopsys translate_off
defparam \Add3~58 .lut_mask = 16'h3C3C;
defparam \Add3~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X55_Y34_N23
dffeas \prif.pc_mem[31] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[31]~2_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[31] .is_wysiwyg = "true";
defparam \prif.pc_mem[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N15
dffeas \prif.rdat1_mem[31] (
	.clk(CLK),
	.d(\PR|rdat1_mem~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[31] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N13
dffeas \prif.pc_bran_mem[31] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [31]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[31] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N8
cycloneive_lcell_comb \Mux101~0 (
// Equation(s):
// \Mux101~0_combout  = (\pc[23]~2_combout  & (((\prif.PCScr_mem [1])))) # (!\pc[23]~2_combout  & ((\prif.PCScr_mem [1] & (\prif.rdat1_mem [31])) # (!\prif.PCScr_mem [1] & ((\prif.pc_bran_mem [31])))))

	.dataa(\pc[23]~2_combout ),
	.datab(\prif.rdat1_mem [31]),
	.datac(\prif.PCScr_mem [1]),
	.datad(\prif.pc_bran_mem [31]),
	.cin(gnd),
	.combout(\Mux101~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux101~0 .lut_mask = 16'hE5E0;
defparam \Mux101~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N6
cycloneive_lcell_comb \Mux101~1 (
// Equation(s):
// \Mux101~1_combout  = (\Mux101~0_combout  & (((\prif.pc_mem [31]) # (!\pc[23]~2_combout )))) # (!\Mux101~0_combout  & (\Add3~58_combout  & ((\pc[23]~2_combout ))))

	.dataa(\Add3~58_combout ),
	.datab(\prif.pc_mem [31]),
	.datac(\Mux101~0_combout ),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux101~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux101~1 .lut_mask = 16'hCAF0;
defparam \Mux101~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X55_Y34_N25
dffeas \prif.pc_mem[30] (
	.clk(CLK),
	.d(\PR|prif.pc_mem[30]~3_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_mem [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_mem[30] .is_wysiwyg = "true";
defparam \prif.pc_mem[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N25
dffeas \prif.pc_bran_mem[30] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[30] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y33_N31
dffeas \prif.rdat1_mem[30] (
	.clk(CLK),
	.d(\PR|rdat1_mem~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [30]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[30] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N10
cycloneive_lcell_comb \Mux102~0 (
// Equation(s):
// \Mux102~0_combout  = (\prif.PCScr_mem [1] & (((\prif.rdat1_mem [30]) # (\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [30] & ((!\pc[23]~2_combout ))))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.pc_bran_mem [30]),
	.datac(\prif.rdat1_mem [30]),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux102~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux102~0 .lut_mask = 16'hAAE4;
defparam \Mux102~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N20
cycloneive_lcell_comb \Mux102~1 (
// Equation(s):
// \Mux102~1_combout  = (\pc[23]~2_combout  & ((\Mux102~0_combout  & (\prif.pc_mem [30])) # (!\Mux102~0_combout  & ((\Add3~56_combout ))))) # (!\pc[23]~2_combout  & (((\Mux102~0_combout ))))

	.dataa(\prif.pc_mem [30]),
	.datab(\Add3~56_combout ),
	.datac(\pc[23]~2_combout ),
	.datad(\Mux102~0_combout ),
	.cin(gnd),
	.combout(\Mux102~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux102~1 .lut_mask = 16'hAFC0;
defparam \Mux102~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y27_N17
dffeas \prif.instr_mem[18] (
	.clk(CLK),
	.d(\PR|instr_mem~17_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[18] .is_wysiwyg = "true";
defparam \prif.instr_mem[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N21
dffeas \prif.rdat1_mem[20] (
	.clk(CLK),
	.d(\PR|rdat1_mem~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [20]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[20] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N18
cycloneive_lcell_comb \Mux112~0 (
// Equation(s):
// \Mux112~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout ) # (\prif.rdat1_mem [20])))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [20] & (!\pc[23]~2_combout )))

	.dataa(\prif.pc_bran_mem [20]),
	.datab(\prif.PCScr_mem [1]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.rdat1_mem [20]),
	.cin(gnd),
	.combout(\Mux112~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux112~0 .lut_mask = 16'hCEC2;
defparam \Mux112~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N24
cycloneive_lcell_comb \Mux112~1 (
// Equation(s):
// \Mux112~1_combout  = (\pc[23]~2_combout  & ((\Mux112~0_combout  & (\prif.instr_mem [18])) # (!\Mux112~0_combout  & ((\Add3~36_combout ))))) # (!\pc[23]~2_combout  & (((\Mux112~0_combout ))))

	.dataa(\prif.instr_mem [18]),
	.datab(\Add3~36_combout ),
	.datac(\pc[23]~2_combout ),
	.datad(\Mux112~0_combout ),
	.cin(gnd),
	.combout(\Mux112~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux112~1 .lut_mask = 16'hAFC0;
defparam \Mux112~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N3
dffeas \prif.pc_bran_mem[17] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[17] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N12
cycloneive_lcell_comb \Mux115~0 (
// Equation(s):
// \Mux115~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & (\Add3~30_combout )) # (!\pc[23]~2_combout  & ((\prif.pc_bran_mem [17])))))

	.dataa(\Add3~30_combout ),
	.datab(\prif.PCScr_mem [1]),
	.datac(\pc[23]~2_combout ),
	.datad(\prif.pc_bran_mem [17]),
	.cin(gnd),
	.combout(\Mux115~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux115~0 .lut_mask = 16'hE3E0;
defparam \Mux115~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N9
dffeas \prif.instr_mem[15] (
	.clk(CLK),
	.d(\PR|instr_mem~18_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [15]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[15] .is_wysiwyg = "true";
defparam \prif.instr_mem[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N5
dffeas \prif.rdat1_mem[17] (
	.clk(CLK),
	.d(\PR|rdat1_mem~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[17] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N10
cycloneive_lcell_comb \Mux115~1 (
// Equation(s):
// \Mux115~1_combout  = (\Mux115~0_combout  & ((\prif.instr_mem [15]) # ((!\prif.PCScr_mem [1])))) # (!\Mux115~0_combout  & (((\prif.rdat1_mem [17] & \prif.PCScr_mem [1]))))

	.dataa(\Mux115~0_combout ),
	.datab(\prif.instr_mem [15]),
	.datac(\prif.rdat1_mem [17]),
	.datad(\prif.PCScr_mem [1]),
	.cin(gnd),
	.combout(\Mux115~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux115~1 .lut_mask = 16'hD8AA;
defparam \Mux115~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y31_N27
dffeas \prif.instr_mem[14] (
	.clk(CLK),
	.d(\PR|instr_mem~19_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [14]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[14] .is_wysiwyg = "true";
defparam \prif.instr_mem[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N15
dffeas \prif.rdat1_mem[16] (
	.clk(CLK),
	.d(\PR|rdat1_mem~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[16] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y31_N29
dffeas \prif.pc_bran_mem[16] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[16] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N6
cycloneive_lcell_comb \Mux116~0 (
// Equation(s):
// \Mux116~0_combout  = (\pc[23]~2_combout  & (\prif.PCScr_mem [1])) # (!\pc[23]~2_combout  & ((\prif.PCScr_mem [1] & (\prif.rdat1_mem [16])) # (!\prif.PCScr_mem [1] & ((\prif.pc_bran_mem [16])))))

	.dataa(\pc[23]~2_combout ),
	.datab(\prif.PCScr_mem [1]),
	.datac(\prif.rdat1_mem [16]),
	.datad(\prif.pc_bran_mem [16]),
	.cin(gnd),
	.combout(\Mux116~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux116~0 .lut_mask = 16'hD9C8;
defparam \Mux116~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N16
cycloneive_lcell_comb \Mux116~1 (
// Equation(s):
// \Mux116~1_combout  = (\pc[23]~2_combout  & ((\Mux116~0_combout  & (\prif.instr_mem [14])) # (!\Mux116~0_combout  & ((\Add3~28_combout ))))) # (!\pc[23]~2_combout  & (((\Mux116~0_combout ))))

	.dataa(\prif.instr_mem [14]),
	.datab(\Add3~28_combout ),
	.datac(\pc[23]~2_combout ),
	.datad(\Mux116~0_combout ),
	.cin(gnd),
	.combout(\Mux116~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux116~1 .lut_mask = 16'hAFC0;
defparam \Mux116~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y30_N11
dffeas \prif.rdat1_mem[19] (
	.clk(CLK),
	.d(\PR|rdat1_mem~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[19] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N1
dffeas \prif.instr_mem[17] (
	.clk(CLK),
	.d(\PR|instr_mem~20_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [17]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[17] .is_wysiwyg = "true";
defparam \prif.instr_mem[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N19
dffeas \prif.pc_bran_mem[19] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~26_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [19]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[19] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N8
cycloneive_lcell_comb \Mux113~0 (
// Equation(s):
// \Mux113~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & (\Add3~34_combout )) # (!\pc[23]~2_combout  & ((\prif.pc_bran_mem [19])))))

	.dataa(\Add3~34_combout ),
	.datab(\prif.pc_bran_mem [19]),
	.datac(\prif.PCScr_mem [1]),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux113~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux113~0 .lut_mask = 16'hFA0C;
defparam \Mux113~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N18
cycloneive_lcell_comb \Mux113~1 (
// Equation(s):
// \Mux113~1_combout  = (\prif.PCScr_mem [1] & ((\Mux113~0_combout  & ((\prif.instr_mem [17]))) # (!\Mux113~0_combout  & (\prif.rdat1_mem [19])))) # (!\prif.PCScr_mem [1] & (((\Mux113~0_combout ))))

	.dataa(\prif.rdat1_mem [19]),
	.datab(\prif.instr_mem [17]),
	.datac(\prif.PCScr_mem [1]),
	.datad(\Mux113~0_combout ),
	.cin(gnd),
	.combout(\Mux113~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux113~1 .lut_mask = 16'hCFA0;
defparam \Mux113~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N9
dffeas \prif.pc_bran_mem[18] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[18] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N3
dffeas \prif.rdat1_mem[18] (
	.clk(CLK),
	.d(\PR|rdat1_mem~27_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [18]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[18] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N22
cycloneive_lcell_comb \Mux114~0 (
// Equation(s):
// \Mux114~0_combout  = (\pc[23]~2_combout  & (\prif.PCScr_mem [1])) # (!\pc[23]~2_combout  & ((\prif.PCScr_mem [1] & ((\prif.rdat1_mem [18]))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [18]))))

	.dataa(\pc[23]~2_combout ),
	.datab(\prif.PCScr_mem [1]),
	.datac(\prif.pc_bran_mem [18]),
	.datad(\prif.rdat1_mem [18]),
	.cin(gnd),
	.combout(\Mux114~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux114~0 .lut_mask = 16'hDC98;
defparam \Mux114~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N11
dffeas \prif.instr_mem[16] (
	.clk(CLK),
	.d(\PR|instr_mem~21_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [16]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[16] .is_wysiwyg = "true";
defparam \prif.instr_mem[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N24
cycloneive_lcell_comb \Mux114~1 (
// Equation(s):
// \Mux114~1_combout  = (\pc[23]~2_combout  & ((\Mux114~0_combout  & (\prif.instr_mem [16])) # (!\Mux114~0_combout  & ((\Add3~32_combout ))))) # (!\pc[23]~2_combout  & (\Mux114~0_combout ))

	.dataa(\pc[23]~2_combout ),
	.datab(\Mux114~0_combout ),
	.datac(\prif.instr_mem [16]),
	.datad(\Add3~32_combout ),
	.cin(gnd),
	.combout(\Mux114~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux114~1 .lut_mask = 16'hE6C4;
defparam \Mux114~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N1
dffeas \prif.rdat1_mem[25] (
	.clk(CLK),
	.d(\PR|rdat1_mem~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[25] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N27
dffeas \prif.pc_bran_mem[25] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~28_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[25] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N14
cycloneive_lcell_comb \Mux107~0 (
// Equation(s):
// \Mux107~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & (\Add3~46_combout )) # (!\pc[23]~2_combout  & ((\prif.pc_bran_mem [25])))))

	.dataa(\Add3~46_combout ),
	.datab(\prif.pc_bran_mem [25]),
	.datac(\prif.PCScr_mem [1]),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux107~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux107~0 .lut_mask = 16'hFA0C;
defparam \Mux107~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N13
dffeas \prif.instr_mem[23] (
	.clk(CLK),
	.d(\PR|instr_mem~22_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [23]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[23] .is_wysiwyg = "true";
defparam \prif.instr_mem[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N4
cycloneive_lcell_comb \Mux107~1 (
// Equation(s):
// \Mux107~1_combout  = (\prif.PCScr_mem [1] & ((\Mux107~0_combout  & ((\prif.instr_mem [23]))) # (!\Mux107~0_combout  & (\prif.rdat1_mem [25])))) # (!\prif.PCScr_mem [1] & (((\Mux107~0_combout ))))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.rdat1_mem [25]),
	.datac(\Mux107~0_combout ),
	.datad(\prif.instr_mem [23]),
	.cin(gnd),
	.combout(\Mux107~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux107~1 .lut_mask = 16'hF858;
defparam \Mux107~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y33_N15
dffeas \prif.instr_mem[22] (
	.clk(CLK),
	.d(\PR|instr_mem~23_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [22]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[22] .is_wysiwyg = "true";
defparam \prif.instr_mem[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N29
dffeas \prif.pc_bran_mem[24] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[24] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X56_Y33_N3
dffeas \prif.rdat1_mem[24] (
	.clk(CLK),
	.d(\PR|rdat1_mem~29_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[24] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N4
cycloneive_lcell_comb \Mux108~0 (
// Equation(s):
// \Mux108~0_combout  = (\prif.PCScr_mem [1] & ((\pc[23]~2_combout ) # ((\prif.rdat1_mem [24])))) # (!\prif.PCScr_mem [1] & (!\pc[23]~2_combout  & (\prif.pc_bran_mem [24])))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\pc[23]~2_combout ),
	.datac(\prif.pc_bran_mem [24]),
	.datad(\prif.rdat1_mem [24]),
	.cin(gnd),
	.combout(\Mux108~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux108~0 .lut_mask = 16'hBA98;
defparam \Mux108~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N30
cycloneive_lcell_comb \Mux108~1 (
// Equation(s):
// \Mux108~1_combout  = (\pc[23]~2_combout  & ((\Mux108~0_combout  & (\prif.instr_mem [22])) # (!\Mux108~0_combout  & ((\Add3~44_combout ))))) # (!\pc[23]~2_combout  & (((\Mux108~0_combout ))))

	.dataa(\prif.instr_mem [22]),
	.datab(\Add3~44_combout ),
	.datac(\pc[23]~2_combout ),
	.datad(\Mux108~0_combout ),
	.cin(gnd),
	.combout(\Mux108~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux108~1 .lut_mask = 16'hAFC0;
defparam \Mux108~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N31
dffeas \prif.instr_mem[25] (
	.clk(CLK),
	.d(\PR|instr_mem~24_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [25]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[25] .is_wysiwyg = "true";
defparam \prif.instr_mem[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y32_N17
dffeas \prif.pc_bran_mem[27] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[27] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N28
cycloneive_lcell_comb \Mux105~0 (
// Equation(s):
// \Mux105~0_combout  = (\prif.PCScr_mem [1] & (((\pc[23]~2_combout )))) # (!\prif.PCScr_mem [1] & ((\pc[23]~2_combout  & ((\Add3~50_combout ))) # (!\pc[23]~2_combout  & (\prif.pc_bran_mem [27]))))

	.dataa(\prif.PCScr_mem [1]),
	.datab(\prif.pc_bran_mem [27]),
	.datac(\Add3~50_combout ),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux105~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux105~0 .lut_mask = 16'hFA44;
defparam \Mux105~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y32_N7
dffeas \prif.rdat1_mem[27] (
	.clk(CLK),
	.d(\PR|rdat1_mem~30_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [27]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[27] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N10
cycloneive_lcell_comb \Mux105~1 (
// Equation(s):
// \Mux105~1_combout  = (\Mux105~0_combout  & ((\prif.instr_mem [25]) # ((!\prif.PCScr_mem [1])))) # (!\Mux105~0_combout  & (((\prif.PCScr_mem [1] & \prif.rdat1_mem [27]))))

	.dataa(\prif.instr_mem [25]),
	.datab(\Mux105~0_combout ),
	.datac(\prif.PCScr_mem [1]),
	.datad(\prif.rdat1_mem [27]),
	.cin(gnd),
	.combout(\Mux105~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux105~1 .lut_mask = 16'hBC8C;
defparam \Mux105~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y32_N25
dffeas \prif.instr_mem[24] (
	.clk(CLK),
	.d(\PR|instr_mem~25_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.instr_mem [24]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.instr_mem[24] .is_wysiwyg = "true";
defparam \prif.instr_mem[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N15
dffeas \prif.pc_bran_mem[26] (
	.clk(CLK),
	.d(\PR|pc_bran_mem~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.pc_bran_mem [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.pc_bran_mem[26] .is_wysiwyg = "true";
defparam \prif.pc_bran_mem[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y32_N29
dffeas \prif.rdat1_mem[26] (
	.clk(CLK),
	.d(\PR|rdat1_mem~31_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.rdat1_mem [26]),
	.prn(vcc));
// synopsys translate_off
defparam \prif.rdat1_mem[26] .is_wysiwyg = "true";
defparam \prif.rdat1_mem[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N16
cycloneive_lcell_comb \Mux106~0 (
// Equation(s):
// \Mux106~0_combout  = (\pc[23]~2_combout  & (\prif.PCScr_mem [1])) # (!\pc[23]~2_combout  & ((\prif.PCScr_mem [1] & ((\prif.rdat1_mem [26]))) # (!\prif.PCScr_mem [1] & (\prif.pc_bran_mem [26]))))

	.dataa(\pc[23]~2_combout ),
	.datab(\prif.PCScr_mem [1]),
	.datac(\prif.pc_bran_mem [26]),
	.datad(\prif.rdat1_mem [26]),
	.cin(gnd),
	.combout(\Mux106~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux106~0 .lut_mask = 16'hDC98;
defparam \Mux106~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N20
cycloneive_lcell_comb \Mux106~1 (
// Equation(s):
// \Mux106~1_combout  = (\Mux106~0_combout  & ((\prif.instr_mem [24]) # ((!\pc[23]~2_combout )))) # (!\Mux106~0_combout  & (((\Add3~48_combout  & \pc[23]~2_combout ))))

	.dataa(\prif.instr_mem [24]),
	.datab(\Mux106~0_combout ),
	.datac(\Add3~48_combout ),
	.datad(\pc[23]~2_combout ),
	.cin(gnd),
	.combout(\Mux106~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux106~1 .lut_mask = 16'hB8CC;
defparam \Mux106~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X52_Y29_N23
dffeas \dpif.halt~_Duplicate_1 (
	.clk(!CLK),
	.d(\dpif.halt~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\dpif.halt~_Duplicate_1_q ),
	.prn(vcc));
// synopsys translate_off
defparam \dpif.halt~_Duplicate_1 .is_wysiwyg = "true";
defparam \dpif.halt~_Duplicate_1 .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y29_N25
dffeas \prif.halt_mem (
	.clk(CLK),
	.d(\PR|halt_mem~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(\prif.rdat1_mem[21]~0_combout ),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\prif.halt_mem~q ),
	.prn(vcc));
// synopsys translate_off
defparam \prif.halt_mem .is_wysiwyg = "true";
defparam \prif.halt_mem .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N22
cycloneive_lcell_comb \dpif.halt~0 (
// Equation(s):
// \dpif.halt~0_combout  = (\dpif.halt~_Duplicate_1_q ) # (\prif.halt_mem~q )

	.dataa(gnd),
	.datab(gnd),
	.datac(\dpif.halt~_Duplicate_1_q ),
	.datad(\prif.halt_mem~q ),
	.cin(gnd),
	.combout(\dpif.halt~0_combout ),
	.cout());
// synopsys translate_off
defparam \dpif.halt~0 .lut_mask = 16'hFFF0;
defparam \dpif.halt~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module alu (
	prifALUOP_ex_3,
	Mux89,
	Mux94,
	Mux30,
	Mux95,
	Mux31,
	Mux92,
	Mux93,
	Mux61,
	Mux91,
	Mux64,
	Mux65,
	Mux66,
	Mux68,
	Mux72,
	Mux77,
	Mux71,
	Mux79,
	Mux76,
	Mux78,
	Mux74,
	Mux75,
	Mux67,
	Mux69,
	Mux73,
	Mux70,
	prifALUOP_ex_2,
	prifALUOP_ex_1,
	Mux29,
	Mux27,
	Mux28,
	Mux931,
	Mux23,
	Mux24,
	Mux25,
	Mux26,
	Mux15,
	Mux16,
	Mux17,
	Mux18,
	Mux20,
	Mux19,
	Mux191,
	Mux21,
	Mux22,
	Mux13,
	Mux14,
	Mux11,
	Mux12,
	Mux9,
	Mux10,
	Mux7,
	Mux8,
	Mux0,
	Mux1,
	Mux2,
	Mux5,
	Mux6,
	Mux3,
	Mux4,
	prifALUOP_ex_0,
	aluifportOut_1,
	Mux192,
	aluifportOut_0,
	aluifportOut_3,
	aluifportOut_5,
	aluifportOut_2,
	aluifportOut_31,
	aluifportOut_32,
	aluifportOut_21,
	aluifportOut_51,
	aluifportOut_52,
	aluifportOut_4,
	aluifportOut_7,
	aluifportOut_6,
	aluifportOut_9,
	aluifportOut_8,
	aluifportOut_11,
	aluifportOut_10,
	aluifportOut_13,
	aluifportOut_12,
	aluifportOut_15,
	aluifportOut_14,
	aluifportOut_23,
	aluifportOut_22,
	aluifportOut_211,
	aluifportOut_29,
	aluifportOut_28,
	aluifneg_flag,
	aluifportOut_30,
	aluifportOut_20,
	aluifportOut_17,
	aluifportOut_16,
	aluifportOut_19,
	aluifportOut_18,
	aluifportOut_25,
	aluifportOut_24,
	aluifportOut_27,
	aluifportOut_26,
	aluifportOut_53,
	Mux90,
	Mux80,
	Mux81,
	Mux82,
	Mux83,
	Mux84,
	Mux85,
	Mux86,
	Mux891,
	Mux87,
	Mux88,
	devpor,
	devclrn,
	devoe);
input 	prifALUOP_ex_3;
input 	Mux89;
input 	Mux94;
input 	Mux30;
input 	Mux95;
input 	Mux31;
input 	Mux92;
input 	Mux93;
input 	Mux61;
input 	Mux91;
input 	Mux64;
input 	Mux65;
input 	Mux66;
input 	Mux68;
input 	Mux72;
input 	Mux77;
input 	Mux71;
input 	Mux79;
input 	Mux76;
input 	Mux78;
input 	Mux74;
input 	Mux75;
input 	Mux67;
input 	Mux69;
input 	Mux73;
input 	Mux70;
input 	prifALUOP_ex_2;
input 	prifALUOP_ex_1;
input 	Mux29;
input 	Mux27;
input 	Mux28;
input 	Mux931;
input 	Mux23;
input 	Mux24;
input 	Mux25;
input 	Mux26;
input 	Mux15;
input 	Mux16;
input 	Mux17;
input 	Mux18;
input 	Mux20;
input 	Mux19;
input 	Mux191;
input 	Mux21;
input 	Mux22;
input 	Mux13;
input 	Mux14;
input 	Mux11;
input 	Mux12;
input 	Mux9;
input 	Mux10;
input 	Mux7;
input 	Mux8;
input 	Mux0;
input 	Mux1;
input 	Mux2;
input 	Mux5;
input 	Mux6;
input 	Mux3;
input 	Mux4;
input 	prifALUOP_ex_0;
output 	aluifportOut_1;
input 	Mux192;
output 	aluifportOut_0;
output 	aluifportOut_3;
output 	aluifportOut_5;
output 	aluifportOut_2;
output 	aluifportOut_31;
output 	aluifportOut_32;
output 	aluifportOut_21;
output 	aluifportOut_51;
output 	aluifportOut_52;
output 	aluifportOut_4;
output 	aluifportOut_7;
output 	aluifportOut_6;
output 	aluifportOut_9;
output 	aluifportOut_8;
output 	aluifportOut_11;
output 	aluifportOut_10;
output 	aluifportOut_13;
output 	aluifportOut_12;
output 	aluifportOut_15;
output 	aluifportOut_14;
output 	aluifportOut_23;
output 	aluifportOut_22;
output 	aluifportOut_211;
output 	aluifportOut_29;
output 	aluifportOut_28;
output 	aluifneg_flag;
output 	aluifportOut_30;
output 	aluifportOut_20;
output 	aluifportOut_17;
output 	aluifportOut_16;
output 	aluifportOut_19;
output 	aluifportOut_18;
output 	aluifportOut_25;
output 	aluifportOut_24;
output 	aluifportOut_27;
output 	aluifportOut_26;
output 	aluifportOut_53;
input 	Mux90;
input 	Mux80;
input 	Mux81;
input 	Mux82;
input 	Mux83;
input 	Mux84;
input 	Mux85;
input 	Mux86;
input 	Mux891;
input 	Mux87;
input 	Mux88;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add0~0_combout ;
wire \Add0~22_combout ;
wire \Add0~26_combout ;
wire \Add0~56_combout ;
wire \ShiftLeft0~8_combout ;
wire \ShiftLeft0~12_combout ;
wire \ShiftRight0~11_combout ;
wire \ShiftRight0~21_combout ;
wire \ShiftRight0~37_combout ;
wire \ShiftRight0~41_combout ;
wire \ShiftRight0~46_combout ;
wire \portOut~0_combout ;
wire \aluif.portOut[0]~19_combout ;
wire \portOut~5_combout ;
wire \portOut~6_combout ;
wire \ShiftRight0~78_combout ;
wire \ShiftRight0~79_combout ;
wire \ShiftRight0~89_combout ;
wire \portOut~9_combout ;
wire \aluif.portOut[5]~53_combout ;
wire \ShiftLeft0~27_combout ;
wire \ShiftLeft0~29_combout ;
wire \ShiftRight0~96_combout ;
wire \portOut~15_combout ;
wire \aluif.portOut[9]~84_combout ;
wire \portOut~25_combout ;
wire \portOut~28_combout ;
wire \ShiftLeft0~52_combout ;
wire \portOut~31_combout ;
wire \aluif.portOut[10]~105_combout ;
wire \portOut~34_combout ;
wire \ShiftLeft0~61_combout ;
wire \portOut~37_combout ;
wire \ShiftRight0~111_combout ;
wire \aluif.portOut[14]~127_combout ;
wire \portOut~42_combout ;
wire \ShiftLeft0~78_combout ;
wire \aluif.portOut[29]~157_combout ;
wire \ShiftLeft0~95_combout ;
wire \aluif.portOut[28]~173_combout ;
wire \aluif.portOut[28]~175_combout ;
wire \portOut~55_combout ;
wire \portOut~56_combout ;
wire \aluif.neg_flag~13_combout ;
wire \aluif.portOut[30]~184_combout ;
wire \aluif.portOut[30]~185_combout ;
wire \portOut~58_combout ;
wire \aluif.portOut[20]~192_combout ;
wire \ShiftLeft0~108_combout ;
wire \aluif.portOut[18]~216_combout ;
wire \aluif.portOut[18]~217_combout ;
wire \aluif.portOut[27]~242_combout ;
wire \aluif.portOut[27]~243_combout ;
wire \aluif.neg_flag~23_combout ;
wire \aluif.portOut[1]~9_combout ;
wire \ShiftLeft0~9_combout ;
wire \ShiftLeft0~11_combout ;
wire \ShiftLeft0~10_combout ;
wire \ShiftLeft0~13_combout ;
wire \ShiftLeft0~14_combout ;
wire \ShiftLeft0~7_combout ;
wire \ShiftLeft0~15_combout ;
wire \ShiftLeft0~5_combout ;
wire \ShiftLeft0~4_combout ;
wire \ShiftLeft0~6_combout ;
wire \aluif.portOut[1]~8_combout ;
wire \Add0~1 ;
wire \Add0~2_combout ;
wire \aluif.portOut[1]~10_combout ;
wire \ShiftRight0~6_combout ;
wire \ShiftRight0~8_combout ;
wire \ShiftRight0~12_combout ;
wire \ShiftRight0~20_combout ;
wire \ShiftRight0~26_combout ;
wire \ShiftLeft0~16_combout ;
wire \ShiftRight0~27_combout ;
wire \ShiftRight0~22_combout ;
wire \ShiftRight0~23_combout ;
wire \ShiftRight0~25_combout ;
wire \ShiftRight0~28_combout ;
wire \ShiftRight0~29_combout ;
wire \ShiftRight0~30_combout ;
wire \ShiftRight0~31_combout ;
wire \ShiftRight0~32_combout ;
wire \aluif.portOut[1]~13_combout ;
wire \Add1~1 ;
wire \Add1~2_combout ;
wire \aluif.portOut[1]~11_combout ;
wire \aluif.portOut[1]~12_combout ;
wire \aluif.portOut[1]~14_combout ;
wire \Add1~0_combout ;
wire \aluif.portOut[0]~16_combout ;
wire \aluif.portOut[0]~17_combout ;
wire \ShiftRight0~53_combout ;
wire \ShiftRight0~54_combout ;
wire \ShiftRight0~55_combout ;
wire \ShiftRight0~57_combout ;
wire \ShiftRight0~56_combout ;
wire \ShiftRight0~58_combout ;
wire \ShiftRight0~59_combout ;
wire \ShiftRight0~50_combout ;
wire \ShiftRight0~49_combout ;
wire \ShiftRight0~51_combout ;
wire \ShiftRight0~47_combout ;
wire \ShiftRight0~48_combout ;
wire \ShiftRight0~52_combout ;
wire \ShiftRight0~60_combout ;
wire \aluif.portOut[0]~18_combout ;
wire \portOut~1_combout ;
wire \aluif.portOut[0]~20_combout ;
wire \aluif.portOut[0]~21_combout ;
wire \aluif.portOut[0]~22_combout ;
wire \LessThan0~1_cout ;
wire \LessThan0~3_cout ;
wire \LessThan0~5_cout ;
wire \LessThan0~7_cout ;
wire \LessThan0~9_cout ;
wire \LessThan0~11_cout ;
wire \LessThan0~13_cout ;
wire \LessThan0~15_cout ;
wire \LessThan0~17_cout ;
wire \LessThan0~19_cout ;
wire \LessThan0~21_cout ;
wire \LessThan0~23_cout ;
wire \LessThan0~25_cout ;
wire \LessThan0~27_cout ;
wire \LessThan0~29_cout ;
wire \LessThan0~31_cout ;
wire \LessThan0~33_cout ;
wire \LessThan0~35_cout ;
wire \LessThan0~37_cout ;
wire \LessThan0~39_cout ;
wire \LessThan0~41_cout ;
wire \LessThan0~43_cout ;
wire \LessThan0~45_cout ;
wire \LessThan0~47_cout ;
wire \LessThan0~49_cout ;
wire \LessThan0~51_cout ;
wire \LessThan0~53_cout ;
wire \LessThan0~55_cout ;
wire \LessThan0~57_cout ;
wire \LessThan0~59_cout ;
wire \LessThan0~61_cout ;
wire \LessThan0~62_combout ;
wire \LessThan1~1_cout ;
wire \LessThan1~3_cout ;
wire \LessThan1~5_cout ;
wire \LessThan1~7_cout ;
wire \LessThan1~9_cout ;
wire \LessThan1~11_cout ;
wire \LessThan1~13_cout ;
wire \LessThan1~15_cout ;
wire \LessThan1~17_cout ;
wire \LessThan1~19_cout ;
wire \LessThan1~21_cout ;
wire \LessThan1~23_cout ;
wire \LessThan1~25_cout ;
wire \LessThan1~27_cout ;
wire \LessThan1~29_cout ;
wire \LessThan1~31_cout ;
wire \LessThan1~33_cout ;
wire \LessThan1~35_cout ;
wire \LessThan1~37_cout ;
wire \LessThan1~39_cout ;
wire \LessThan1~41_cout ;
wire \LessThan1~43_cout ;
wire \LessThan1~45_cout ;
wire \LessThan1~47_cout ;
wire \LessThan1~49_cout ;
wire \LessThan1~51_cout ;
wire \LessThan1~53_cout ;
wire \LessThan1~55_cout ;
wire \LessThan1~57_cout ;
wire \LessThan1~59_cout ;
wire \LessThan1~61_cout ;
wire \LessThan1~62_combout ;
wire \aluif.portOut[0]~23_combout ;
wire \portOut~4_combout ;
wire \aluif.portOut[5]~25_combout ;
wire \aluif.portOut[2]~29_combout ;
wire \Add0~3 ;
wire \Add0~5 ;
wire \Add0~6_combout ;
wire \portOut~2_combout ;
wire \aluif.portOut[15]~26_combout ;
wire \portOut~3_combout ;
wire \aluif.portOut[3]~27_combout ;
wire \aluif.portOut[3]~28_combout ;
wire \aluif.portOut[2]~32_combout ;
wire \Add1~3 ;
wire \Add1~5 ;
wire \Add1~6_combout ;
wire \aluif.portOut[2]~34_combout ;
wire \aluif.portOut[2]~35_combout ;
wire \ShiftRight0~10_combout ;
wire \ShiftRight0~61_combout ;
wire \ShiftRight0~17_combout ;
wire \ShiftRight0~9_combout ;
wire \ShiftRight0~72_combout ;
wire \ShiftRight0~7_combout ;
wire \aluif.portOut[3]~36_combout ;
wire \aluif.portOut[3]~37_combout ;
wire \ShiftRight0~62_combout ;
wire \ShiftRight0~63_combout ;
wire \ShiftRight0~65_combout ;
wire \ShiftRight0~66_combout ;
wire \ShiftRight0~67_combout ;
wire \ShiftRight0~70_combout ;
wire \ShiftRight0~71_combout ;
wire \aluif.portOut[3]~38_combout ;
wire \Add1~4_combout ;
wire \ShiftRight0~90_combout ;
wire \ShiftRight0~88_combout ;
wire \ShiftRight0~91_combout ;
wire \ShiftRight0~87_combout ;
wire \aluif.portOut[2]~44_combout ;
wire \aluif.portOut[2]~45_combout ;
wire \portOut~7_combout ;
wire \aluif.portOut[2]~46_combout ;
wire \ShiftRight0~77_combout ;
wire \ShiftRight0~80_combout ;
wire \ShiftRight0~81_combout ;
wire \ShiftRight0~82_combout ;
wire \ShiftRight0~85_combout ;
wire \ShiftRight0~86_combout ;
wire \aluif.portOut[2]~47_combout ;
wire \Add0~4_combout ;
wire \ShiftLeft0~20_combout ;
wire \ShiftLeft0~21_combout ;
wire \ShiftLeft0~109_combout ;
wire \aluif.portOut[2]~41_combout ;
wire \aluif.portOut[2]~42_combout ;
wire \aluif.portOut[2]~43_combout ;
wire \Add1~7 ;
wire \Add1~9 ;
wire \Add1~10_combout ;
wire \portOut~10_combout ;
wire \aluif.portOut[5]~55_combout ;
wire \aluif.portOut[5]~51_combout ;
wire \ShiftRight0~93_combout ;
wire \ShiftRight0~24_combout ;
wire \ShiftRight0~94_combout ;
wire \ShiftRight0~112_combout ;
wire \ShiftRight0~95_combout ;
wire \ShiftRight0~14_combout ;
wire \ShiftRight0~13_combout ;
wire \ShiftRight0~15_combout ;
wire \ShiftRight0~92_combout ;
wire \aluif.portOut[5]~54_combout ;
wire \aluif.portOut[5]~56_combout ;
wire \Add0~7 ;
wire \Add0~9 ;
wire \Add0~10_combout ;
wire \ShiftLeft0~18_combout ;
wire \ShiftLeft0~23_combout ;
wire \ShiftLeft0~24_combout ;
wire \ShiftLeft0~22_combout ;
wire \ShiftLeft0~25_combout ;
wire \aluif.portOut[5]~49_combout ;
wire \portOut~8_combout ;
wire \aluif.portOut[5]~50_combout ;
wire \Add0~8_combout ;
wire \portOut~11_combout ;
wire \portOut~12_combout ;
wire \aluif.portOut[4]~59_combout ;
wire \aluif.portOut[4]~60_combout ;
wire \portOut~13_combout ;
wire \Add1~8_combout ;
wire \aluif.portOut[5]~52_combout ;
wire \aluif.portOut[4]~61_combout ;
wire \ShiftRight0~43_combout ;
wire \ShiftRight0~44_combout ;
wire \ShiftRight0~98_combout ;
wire \aluif.portOut[4]~62_combout ;
wire \aluif.portOut[4]~63_combout ;
wire \aluif.portOut[4]~64_combout ;
wire \ShiftRight0~75_combout ;
wire \ShiftRight0~74_combout ;
wire \ShiftRight0~68_combout ;
wire \ShiftRight0~69_combout ;
wire \ShiftRight0~99_combout ;
wire \aluif.portOut[7]~68_combout ;
wire \ShiftRight0~16_combout ;
wire \ShiftRight0~73_combout ;
wire \ShiftRight0~64_combout ;
wire \ShiftRight0~100_combout ;
wire \ShiftRight0~101_combout ;
wire \aluif.portOut[7]~69_combout ;
wire \aluif.portOut[7]~70_combout ;
wire \Add1~11 ;
wire \Add1~13 ;
wire \Add1~14_combout ;
wire \portOut~16_combout ;
wire \aluif.portOut[7]~71_combout ;
wire \Add0~11 ;
wire \Add0~13 ;
wire \Add0~14_combout ;
wire \portOut~14_combout ;
wire \ShiftLeft0~31_combout ;
wire \ShiftLeft0~32_combout ;
wire \ShiftLeft0~30_combout ;
wire \ShiftLeft0~33_combout ;
wire \aluif.portOut[7]~66_combout ;
wire \aluif.portOut[7]~67_combout ;
wire \Add0~12_combout ;
wire \portOut~17_combout ;
wire \ShiftLeft0~34_combout ;
wire \ShiftLeft0~35_combout ;
wire \ShiftLeft0~36_combout ;
wire \portOut~18_combout ;
wire \aluif.portOut[6]~73_combout ;
wire \aluif.portOut[6]~74_combout ;
wire \Add1~12_combout ;
wire \portOut~19_combout ;
wire \ShiftRight0~103_combout ;
wire \ShiftRight0~104_combout ;
wire \ShiftRight0~83_combout ;
wire \ShiftRight0~84_combout ;
wire \ShiftRight0~102_combout ;
wire \aluif.portOut[6]~75_combout ;
wire \aluif.portOut[6]~76_combout ;
wire \aluif.portOut[6]~77_combout ;
wire \aluif.portOut[6]~78_combout ;
wire \Add1~15 ;
wire \Add1~17 ;
wire \Add1~18_combout ;
wire \aluif.portOut[15]~80_combout ;
wire \ShiftRight0~18_combout ;
wire \ShiftRight0~19_combout ;
wire \aluif.portOut[15]~81_combout ;
wire \aluif.portOut[9]~85_combout ;
wire \aluif.portOut[15]~86_combout ;
wire \portOut~21_combout ;
wire \Add0~15 ;
wire \Add0~17 ;
wire \Add0~18_combout ;
wire \portOut~22_combout ;
wire \ShiftLeft0~37_combout ;
wire \ShiftLeft0~38_combout ;
wire \ShiftLeft0~39_combout ;
wire \ShiftLeft0~40_combout ;
wire \aluif.portOut[9]~87_combout ;
wire \aluif.portOut[9]~88_combout ;
wire \aluif.portOut[9]~89_combout ;
wire \portOut~20_combout ;
wire \portOut~23_combout ;
wire \Add1~16_combout ;
wire \portOut~24_combout ;
wire \Add0~16_combout ;
wire \ShiftLeft0~110_combout ;
wire \ShiftLeft0~26_combout ;
wire \ShiftLeft0~28_combout ;
wire \ShiftLeft0~41_combout ;
wire \ShiftLeft0~42_combout ;
wire \ShiftLeft0~43_combout ;
wire \ShiftLeft0~44_combout ;
wire \aluif.portOut[8]~93_combout ;
wire \aluif.portOut[8]~94_combout ;
wire \aluif.portOut[8]~95_combout ;
wire \ShiftRight0~36_combout ;
wire \ShiftRight0~34_combout ;
wire \ShiftRight0~33_combout ;
wire \ShiftRight0~35_combout ;
wire \ShiftRight0~38_combout ;
wire \ShiftRight0~106_combout ;
wire \aluif.portOut[15]~82_combout ;
wire \aluif.portOut[15]~83_combout ;
wire \aluif.portOut[8]~91_combout ;
wire \aluif.portOut[8]~92_combout ;
wire \portOut~26_combout ;
wire \ShiftRight0~76_combout ;
wire \ShiftRight0~107_combout ;
wire \aluif.portOut[11]~97_combout ;
wire \aluif.portOut[11]~98_combout ;
wire \portOut~27_combout ;
wire \ShiftLeft0~46_combout ;
wire \ShiftLeft0~47_combout ;
wire \ShiftLeft0~48_combout ;
wire \aluif.portOut[11]~99_combout ;
wire \aluif.portOut[11]~100_combout ;
wire \aluif.portOut[11]~101_combout ;
wire \Add1~19 ;
wire \Add1~21 ;
wire \Add1~22_combout ;
wire \portOut~29_combout ;
wire \Add1~20_combout ;
wire \portOut~30_combout ;
wire \Add0~19 ;
wire \Add0~20_combout ;
wire \aluif.portOut[10]~106_combout ;
wire \aluif.portOut[10]~107_combout ;
wire \ShiftRight0~108_combout ;
wire \aluif.portOut[10]~103_combout ;
wire \aluif.portOut[10]~104_combout ;
wire \ShiftRight0~109_combout ;
wire \portOut~32_combout ;
wire \aluif.portOut[13]~109_combout ;
wire \aluif.portOut[13]~110_combout ;
wire \portOut~33_combout ;
wire \ShiftLeft0~53_combout ;
wire \ShiftLeft0~45_combout ;
wire \ShiftLeft0~55_combout ;
wire \ShiftLeft0~56_combout ;
wire \ShiftLeft0~57_combout ;
wire \aluif.portOut[13]~111_combout ;
wire \aluif.portOut[13]~112_combout ;
wire \Add1~23 ;
wire \Add1~25 ;
wire \Add1~26_combout ;
wire \aluif.portOut[13]~113_combout ;
wire \Add1~24_combout ;
wire \portOut~35_combout ;
wire \Add0~21 ;
wire \Add0~23 ;
wire \Add0~24_combout ;
wire \ShiftLeft0~58_combout ;
wire \ShiftLeft0~62_combout ;
wire \aluif.portOut[12]~117_combout ;
wire \portOut~36_combout ;
wire \aluif.portOut[12]~118_combout ;
wire \ShiftRight0~39_combout ;
wire \ShiftRight0~40_combout ;
wire \ShiftRight0~97_combout ;
wire \ShiftRight0~42_combout ;
wire \ShiftRight0~110_combout ;
wire \aluif.portOut[12]~115_combout ;
wire \aluif.portOut[12]~116_combout ;
wire \aluif.portOut[12]~119_combout ;
wire \portOut~38_combout ;
wire \Add1~27 ;
wire \Add1~29 ;
wire \Add1~30_combout ;
wire \portOut~39_combout ;
wire \Add0~25 ;
wire \Add0~27 ;
wire \Add0~29 ;
wire \Add0~30_combout ;
wire \ShiftLeft0~63_combout ;
wire \ShiftLeft0~54_combout ;
wire \ShiftLeft0~64_combout ;
wire \ShiftLeft0~65_combout ;
wire \ShiftLeft0~66_combout ;
wire \ShiftLeft0~67_combout ;
wire \portOut~40_combout ;
wire \aluif.portOut[15]~123_combout ;
wire \aluif.portOut[15]~124_combout ;
wire \aluif.portOut[15]~125_combout ;
wire \ShiftRight0~113_combout ;
wire \aluif.portOut[15]~121_combout ;
wire \aluif.portOut[15]~122_combout ;
wire \Add1~28_combout ;
wire \portOut~41_combout ;
wire \Add0~28_combout ;
wire \portOut~43_combout ;
wire \aluif.portOut[14]~129_combout ;
wire \aluif.portOut[14]~130_combout ;
wire \aluif.portOut[14]~128_combout ;
wire \aluif.portOut[14]~131_combout ;
wire \Add1~31 ;
wire \Add1~33 ;
wire \Add1~35 ;
wire \Add1~37 ;
wire \Add1~39 ;
wire \Add1~41 ;
wire \Add1~43 ;
wire \Add1~45 ;
wire \Add1~46_combout ;
wire \portOut~44_combout ;
wire \aluif.portOut[23]~133_combout ;
wire \aluif.portOut[23]~134_combout ;
wire \portOut~46_combout ;
wire \aluif.portOut[23]~135_combout ;
wire \aluif.portOut[23]~136_combout ;
wire \ShiftLeft0~75_combout ;
wire \ShiftLeft0~73_combout ;
wire \ShiftLeft0~74_combout ;
wire \ShiftLeft0~77_combout ;
wire \portOut~45_combout ;
wire \aluif.portOut[23]~137_combout ;
wire \aluif.portOut[23]~138_combout ;
wire \Add0~31 ;
wire \Add0~33 ;
wire \Add0~35 ;
wire \Add0~37 ;
wire \Add0~39 ;
wire \Add0~41 ;
wire \Add0~43 ;
wire \Add0~45 ;
wire \Add0~46_combout ;
wire \aluif.portOut[23]~139_combout ;
wire \aluif.portOut[22]~144_combout ;
wire \portOut~48_combout ;
wire \aluif.portOut[22]~143_combout ;
wire \aluif.portOut[22]~259_combout ;
wire \ShiftLeft0~49_combout ;
wire \ShiftLeft0~50_combout ;
wire \ShiftLeft0~59_combout ;
wire \ShiftLeft0~69_combout ;
wire \ShiftLeft0~70_combout ;
wire \ShiftLeft0~71_combout ;
wire \portOut~47_combout ;
wire \aluif.portOut[22]~141_combout ;
wire \ShiftLeft0~80_combout ;
wire \ShiftLeft0~79_combout ;
wire \ShiftLeft0~81_combout ;
wire \ShiftLeft0~82_combout ;
wire \aluif.portOut[22]~142_combout ;
wire \aluif.portOut[22]~145_combout ;
wire \Add0~44_combout ;
wire \Add1~44_combout ;
wire \aluif.portOut[22]~260_combout ;
wire \aluif.portOut[22]~146_combout ;
wire \aluif.portOut[22]~261_combout ;
wire \portOut~51_combout ;
wire \portOut~49_combout ;
wire \Add1~42_combout ;
wire \aluif.portOut[21]~148_combout ;
wire \aluif.portOut[21]~149_combout ;
wire \Add0~42_combout ;
wire \ShiftLeft0~83_combout ;
wire \ShiftLeft0~84_combout ;
wire \ShiftLeft0~85_combout ;
wire \ShiftLeft0~86_combout ;
wire \ShiftLeft0~87_combout ;
wire \portOut~50_combout ;
wire \aluif.portOut[21]~150_combout ;
wire \aluif.portOut[21]~151_combout ;
wire \aluif.portOut[21]~152_combout ;
wire \aluif.portOut[28]~154_combout ;
wire \Add1~47 ;
wire \Add1~49 ;
wire \Add1~51 ;
wire \Add1~53 ;
wire \Add1~55 ;
wire \Add1~57 ;
wire \Add1~58_combout ;
wire \aluif.portOut[29]~164_combout ;
wire \portOut~52_combout ;
wire \aluif.portOut[29]~155_combout ;
wire \aluif.portOut[29]~163_combout ;
wire \aluif.portOut[29]~165_combout ;
wire \ShiftLeft0~88_combout ;
wire \aluif.portOut[29]~158_combout ;
wire \aluif.portOut[29]~159_combout ;
wire \Add0~47 ;
wire \Add0~49 ;
wire \Add0~51 ;
wire \Add0~53 ;
wire \Add0~55 ;
wire \Add0~57 ;
wire \Add0~58_combout ;
wire \aluif.portOut[29]~160_combout ;
wire \aluif.portOut[29]~162_combout ;
wire \aluif.portOut[29]~156_combout ;
wire \aluif.portOut[29]~161_combout ;
wire \aluif.portOut[28]~168_combout ;
wire \aluif.portOut[28]~171_combout ;
wire \aluif.portOut[28]~262_combout ;
wire \ShiftLeft0~92_combout ;
wire \ShiftLeft0~96_combout ;
wire \ShiftLeft0~97_combout ;
wire \ShiftLeft0~99_combout ;
wire \ShiftLeft0~100_combout ;
wire \aluif.portOut[28]~174_combout ;
wire \aluif.portOut[28]~177_combout ;
wire \portOut~53_combout ;
wire \aluif.portOut[28]~172_combout ;
wire \aluif.portOut[28]~176_combout ;
wire \aluif.portOut[28]~178_combout ;
wire \aluif.portOut[28]~169_combout ;
wire \aluif.portOut[28]~170_combout ;
wire \aluif.portOut[28]~179_combout ;
wire \aluif.portOut[28]~167_combout ;
wire \Add1~56_combout ;
wire \Add0~59 ;
wire \Add0~61 ;
wire \Add0~62_combout ;
wire \Add1~59 ;
wire \Add1~61 ;
wire \Add1~62_combout ;
wire \portOut~54_combout ;
wire \aluif.neg_flag~12_combout ;
wire \aluif.neg_flag~21_combout ;
wire \ShiftLeft0~101_combout ;
wire \ShiftLeft0~102_combout ;
wire \aluif.portOut[30]~181_combout ;
wire \ShiftLeft0~91_combout ;
wire \aluif.neg_flag~14_combout ;
wire \aluif.neg_flag~15_combout ;
wire \aluif.neg_flag~16_combout ;
wire \aluif.neg_flag~18_combout ;
wire \aluif.neg_flag~20_combout ;
wire \aluif.neg_flag~17_combout ;
wire \aluif.neg_flag~22_combout ;
wire \portOut~59_combout ;
wire \Add1~60_combout ;
wire \portOut~57_combout ;
wire \aluif.portOut[30]~182_combout ;
wire \aluif.portOut[30]~183_combout ;
wire \Add0~60_combout ;
wire \ShiftLeft0~68_combout ;
wire \ShiftLeft0~72_combout ;
wire \aluif.portOut[30]~186_combout ;
wire \aluif.portOut[30]~187_combout ;
wire \aluif.portOut[30]~188_combout ;
wire \portOut~62_combout ;
wire \Add0~40_combout ;
wire \portOut~60_combout ;
wire \aluif.portOut[20]~190_combout ;
wire \aluif.portOut[20]~191_combout ;
wire \Add1~40_combout ;
wire \portOut~61_combout ;
wire \aluif.portOut[20]~193_combout ;
wire \aluif.portOut[20]~194_combout ;
wire \Add0~34_combout ;
wire \portOut~65_combout ;
wire \portOut~63_combout ;
wire \aluif.portOut[17]~196_combout ;
wire \Add1~34_combout ;
wire \aluif.portOut[17]~197_combout ;
wire \portOut~64_combout ;
wire \aluif.portOut[17]~198_combout ;
wire \ShiftLeft0~105_combout ;
wire \aluif.portOut[17]~199_combout ;
wire \aluif.portOut[17]~200_combout ;
wire \Add0~32_combout ;
wire \ShiftLeft0~98_combout ;
wire \ShiftLeft0~60_combout ;
wire \ShiftLeft0~106_combout ;
wire \ShiftLeft0~17_combout ;
wire \portOut~67_combout ;
wire \aluif.portOut[16]~204_combout ;
wire \aluif.portOut[16]~205_combout ;
wire \aluif.portOut[16]~206_combout ;
wire \portOut~68_combout ;
wire \portOut~66_combout ;
wire \ShiftRight0~45_combout ;
wire \aluif.portOut[16]~202_combout ;
wire \Add1~32_combout ;
wire \aluif.portOut[16]~203_combout ;
wire \portOut~71_combout ;
wire \ShiftLeft0~76_combout ;
wire \ShiftLeft0~107_combout ;
wire \ShiftLeft0~19_combout ;
wire \portOut~70_combout ;
wire \aluif.portOut[19]~210_combout ;
wire \aluif.portOut[19]~211_combout ;
wire \Add0~38_combout ;
wire \aluif.portOut[19]~212_combout ;
wire \Add1~38_combout ;
wire \portOut~69_combout ;
wire \aluif.portOut[19]~208_combout ;
wire \aluif.portOut[19]~209_combout ;
wire \portOut~74_combout ;
wire \Add0~36_combout ;
wire \portOut~73_combout ;
wire \aluif.portOut[18]~218_combout ;
wire \ShiftLeft0~51_combout ;
wire \aluif.portOut[18]~219_combout ;
wire \portOut~72_combout ;
wire \Add1~36_combout ;
wire \aluif.portOut[18]~214_combout ;
wire \aluif.portOut[18]~215_combout ;
wire \aluif.portOut[18]~220_combout ;
wire \aluif.portOut[25]~226_combout ;
wire \ShiftLeft0~89_combout ;
wire \ShiftLeft0~90_combout ;
wire \aluif.portOut[25]~222_combout ;
wire \aluif.portOut[25]~223_combout ;
wire \ShiftRight0~105_combout ;
wire \aluif.portOut[25]~227_combout ;
wire \aluif.portOut[25]~228_combout ;
wire \aluif.portOut[25]~229_combout ;
wire \aluif.portOut[25]~225_combout ;
wire \aluif.portOut[25]~230_combout ;
wire \aluif.portOut[25]~231_combout ;
wire \aluif.portOut[25]~232_combout ;
wire \Add1~50_combout ;
wire \aluif.portOut[25]~233_combout ;
wire \Add0~50_combout ;
wire \portOut~75_combout ;
wire \aluif.portOut[25]~224_combout ;
wire \portOut~77_combout ;
wire \ShiftLeft0~93_combout ;
wire \ShiftLeft0~94_combout ;
wire \aluif.portOut[24]~235_combout ;
wire \aluif.portOut[24]~236_combout ;
wire \aluif.portOut[24]~237_combout ;
wire \Add0~48_combout ;
wire \portOut~76_combout ;
wire \aluif.portOut[24]~238_combout ;
wire \portOut~78_combout ;
wire \Add1~48_combout ;
wire \aluif.portOut[24]~239_combout ;
wire \aluif.portOut[24]~240_combout ;
wire \portOut~80_combout ;
wire \Add1~54_combout ;
wire \aluif.portOut[27]~247_combout ;
wire \aluif.portOut[27]~248_combout ;
wire \Add0~54_combout ;
wire \aluif.portOut[27]~245_combout ;
wire \portOut~79_combout ;
wire \aluif.portOut[27]~244_combout ;
wire \aluif.portOut[27]~246_combout ;
wire \portOut~82_combout ;
wire \Add1~52_combout ;
wire \aluif.portOut[26]~255_combout ;
wire \aluif.portOut[26]~256_combout ;
wire \Add0~52_combout ;
wire \aluif.portOut[26]~253_combout ;
wire \portOut~81_combout ;
wire \ShiftLeft0~103_combout ;
wire \ShiftLeft0~104_combout ;
wire \aluif.portOut[26]~250_combout ;
wire \aluif.portOut[26]~251_combout ;
wire \aluif.portOut[26]~252_combout ;
wire \aluif.portOut[26]~254_combout ;


// Location: LCCOMB_X55_Y25_N0
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = (\Mux31~1_combout  & (\Mux95~1_combout  $ (VCC))) # (!\Mux31~1_combout  & (\Mux95~1_combout  & VCC))
// \Add0~1  = CARRY((\Mux31~1_combout  & \Mux95~1_combout ))

	.dataa(Mux31),
	.datab(Mux95),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout(\Add0~1 ));
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h6688;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N22
cycloneive_lcell_comb \Add0~22 (
// Equation(s):
// \Add0~22_combout  = (\Mux84~3_combout  & ((\Mux20~1_combout  & (\Add0~21  & VCC)) # (!\Mux20~1_combout  & (!\Add0~21 )))) # (!\Mux84~3_combout  & ((\Mux20~1_combout  & (!\Add0~21 )) # (!\Mux20~1_combout  & ((\Add0~21 ) # (GND)))))
// \Add0~23  = CARRY((\Mux84~3_combout  & (!\Mux20~1_combout  & !\Add0~21 )) # (!\Mux84~3_combout  & ((!\Add0~21 ) # (!\Mux20~1_combout ))))

	.dataa(Mux84),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~21 ),
	.combout(\Add0~22_combout ),
	.cout(\Add0~23 ));
// synopsys translate_off
defparam \Add0~22 .lut_mask = 16'h9617;
defparam \Add0~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N26
cycloneive_lcell_comb \Add0~26 (
// Equation(s):
// \Add0~26_combout  = (\Mux82~3_combout  & ((\Mux18~1_combout  & (\Add0~25  & VCC)) # (!\Mux18~1_combout  & (!\Add0~25 )))) # (!\Mux82~3_combout  & ((\Mux18~1_combout  & (!\Add0~25 )) # (!\Mux18~1_combout  & ((\Add0~25 ) # (GND)))))
// \Add0~27  = CARRY((\Mux82~3_combout  & (!\Mux18~1_combout  & !\Add0~25 )) # (!\Mux82~3_combout  & ((!\Add0~25 ) # (!\Mux18~1_combout ))))

	.dataa(Mux82),
	.datab(Mux18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~25 ),
	.combout(\Add0~26_combout ),
	.cout(\Add0~27 ));
// synopsys translate_off
defparam \Add0~26 .lut_mask = 16'h9617;
defparam \Add0~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N24
cycloneive_lcell_comb \Add0~56 (
// Equation(s):
// \Add0~56_combout  = ((\Mux67~0_combout  $ (\Mux3~1_combout  $ (!\Add0~55 )))) # (GND)
// \Add0~57  = CARRY((\Mux67~0_combout  & ((\Mux3~1_combout ) # (!\Add0~55 ))) # (!\Mux67~0_combout  & (\Mux3~1_combout  & !\Add0~55 )))

	.dataa(Mux67),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~55 ),
	.combout(\Add0~56_combout ),
	.cout(\Add0~57 ));
// synopsys translate_off
defparam \Add0~56 .lut_mask = 16'h698E;
defparam \Add0~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N30
cycloneive_lcell_comb \ShiftLeft0~8 (
// Equation(s):
// \ShiftLeft0~8_combout  = (\Mux90~3_combout ) # ((\Mux82~3_combout ) # ((\Mux81~3_combout ) # (\Mux80~4_combout )))

	.dataa(Mux90),
	.datab(Mux82),
	.datac(Mux81),
	.datad(Mux80),
	.cin(gnd),
	.combout(\ShiftLeft0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~8 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N6
cycloneive_lcell_comb \ShiftLeft0~12 (
// Equation(s):
// \ShiftLeft0~12_combout  = (\Mux69~0_combout ) # ((\Mux75~0_combout ) # ((\Mux74~0_combout ) # (\Mux67~0_combout )))

	.dataa(Mux69),
	.datab(Mux75),
	.datac(Mux74),
	.datad(Mux67),
	.cin(gnd),
	.combout(\ShiftLeft0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~12 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N30
cycloneive_lcell_comb \ShiftRight0~11 (
// Equation(s):
// \ShiftRight0~11_combout  = (\Mux94~1_combout  & (\ShiftRight0~9_combout )) # (!\Mux94~1_combout  & ((\ShiftRight0~10_combout )))

	.dataa(Mux94),
	.datab(gnd),
	.datac(\ShiftRight0~9_combout ),
	.datad(\ShiftRight0~10_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~11 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N26
cycloneive_lcell_comb \ShiftRight0~21 (
// Equation(s):
// \ShiftRight0~21_combout  = (\Mux95~1_combout  & ((\Mux11~1_combout ) # ((!\Mux94~1_combout )))) # (!\Mux95~1_combout  & (((\Mux12~1_combout  & \Mux94~1_combout ))))

	.dataa(Mux95),
	.datab(Mux11),
	.datac(Mux12),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftRight0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~21 .lut_mask = 16'hD8AA;
defparam \ShiftRight0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N22
cycloneive_lcell_comb \ShiftRight0~37 (
// Equation(s):
// \ShiftRight0~37_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux8~1_combout ))) # (!\Mux95~1_combout  & (\Mux9~1_combout ))))

	.dataa(Mux94),
	.datab(Mux9),
	.datac(Mux8),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~37 .lut_mask = 16'hA088;
defparam \ShiftRight0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N26
cycloneive_lcell_comb \ShiftRight0~41 (
// Equation(s):
// \ShiftRight0~41_combout  = (\Mux92~2_combout  & (\ShiftRight0~40_combout  & (!\Mux93~2_combout ))) # (!\Mux92~2_combout  & (((\ShiftRight0~38_combout ))))

	.dataa(\ShiftRight0~40_combout ),
	.datab(Mux931),
	.datac(Mux92),
	.datad(\ShiftRight0~38_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~41 .lut_mask = 16'h2F20;
defparam \ShiftRight0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N6
cycloneive_lcell_comb \ShiftRight0~46 (
// Equation(s):
// \ShiftRight0~46_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux30~1_combout ))) # (!\Mux95~1_combout  & (\Mux31~1_combout ))))

	.dataa(Mux94),
	.datab(Mux31),
	.datac(Mux30),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~46 .lut_mask = 16'h5044;
defparam \ShiftRight0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y23_N24
cycloneive_lcell_comb \portOut~0 (
// Equation(s):
// \portOut~0_combout  = (\Mux31~1_combout  & \Mux95~1_combout )

	.dataa(gnd),
	.datab(Mux31),
	.datac(gnd),
	.datad(Mux95),
	.cin(gnd),
	.combout(\portOut~0_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~0 .lut_mask = 16'hCC00;
defparam \portOut~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N12
cycloneive_lcell_comb \aluif.portOut[0]~19 (
// Equation(s):
// \aluif.portOut[0]~19_combout  = (\prif.ALUOP_ex [2] & (!\Mux91~2_combout  & ((\ShiftLeft0~17_combout )))) # (!\prif.ALUOP_ex [2] & (((\portOut~0_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(Mux91),
	.datac(\portOut~0_combout ),
	.datad(\ShiftLeft0~17_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[0]~19_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[0]~19 .lut_mask = 16'h7250;
defparam \aluif.portOut[0]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N30
cycloneive_lcell_comb \portOut~5 (
// Equation(s):
// \portOut~5_combout  = \Mux93~2_combout  $ (\Mux29~1_combout )

	.dataa(gnd),
	.datab(Mux931),
	.datac(Mux29),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~5_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~5 .lut_mask = 16'h3C3C;
defparam \portOut~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N2
cycloneive_lcell_comb \portOut~6 (
// Equation(s):
// \portOut~6_combout  = (\Mux93~2_combout  & \Mux29~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux931),
	.datad(Mux29),
	.cin(gnd),
	.combout(\portOut~6_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~6 .lut_mask = 16'hF000;
defparam \portOut~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N24
cycloneive_lcell_comb \ShiftRight0~78 (
// Equation(s):
// \ShiftRight0~78_combout  = (\Mux95~1_combout  & (\Mux94~1_combout )) # (!\Mux95~1_combout  & ((\Mux94~1_combout  & (\Mux3~1_combout )) # (!\Mux94~1_combout  & ((\Mux5~1_combout )))))

	.dataa(Mux95),
	.datab(Mux94),
	.datac(Mux3),
	.datad(Mux5),
	.cin(gnd),
	.combout(\ShiftRight0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~78 .lut_mask = 16'hD9C8;
defparam \ShiftRight0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N6
cycloneive_lcell_comb \ShiftRight0~79 (
// Equation(s):
// \ShiftRight0~79_combout  = (\ShiftRight0~78_combout  & (((\Mux2~1_combout ) # (!\Mux95~1_combout )))) # (!\ShiftRight0~78_combout  & (\Mux4~1_combout  & ((\Mux95~1_combout ))))

	.dataa(Mux4),
	.datab(\ShiftRight0~78_combout ),
	.datac(Mux2),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~79 .lut_mask = 16'hE2CC;
defparam \ShiftRight0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N26
cycloneive_lcell_comb \ShiftRight0~89 (
// Equation(s):
// \ShiftRight0~89_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux16~1_combout )) # (!\Mux95~1_combout  & ((\Mux17~1_combout )))))

	.dataa(Mux94),
	.datab(Mux95),
	.datac(Mux16),
	.datad(Mux17),
	.cin(gnd),
	.combout(\ShiftRight0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~89 .lut_mask = 16'h5140;
defparam \ShiftRight0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N22
cycloneive_lcell_comb \portOut~9 (
// Equation(s):
// \portOut~9_combout  = (\Mux90~3_combout  & \Mux26~1_combout )

	.dataa(gnd),
	.datab(Mux90),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\portOut~9_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~9 .lut_mask = 16'hCC00;
defparam \portOut~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N6
cycloneive_lcell_comb \aluif.portOut[5]~53 (
// Equation(s):
// \aluif.portOut[5]~53_combout  = (\aluif.portOut[5]~51_combout  & (((\aluif.portOut[5]~52_combout )))) # (!\aluif.portOut[5]~51_combout  & ((\aluif.portOut[5]~52_combout  & ((\ShiftRight0~18_combout ))) # (!\aluif.portOut[5]~52_combout  & 
// (\ShiftRight0~11_combout ))))

	.dataa(\ShiftRight0~11_combout ),
	.datab(\aluif.portOut[5]~51_combout ),
	.datac(\aluif.portOut[5]~52_combout ),
	.datad(\ShiftRight0~18_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[5]~53_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~53 .lut_mask = 16'hF2C2;
defparam \aluif.portOut[5]~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N6
cycloneive_lcell_comb \ShiftLeft0~27 (
// Equation(s):
// \ShiftLeft0~27_combout  = (\Mux95~1_combout  & (\Mux28~1_combout )) # (!\Mux95~1_combout  & ((\Mux27~1_combout )))

	.dataa(Mux28),
	.datab(Mux95),
	.datac(gnd),
	.datad(Mux27),
	.cin(gnd),
	.combout(\ShiftLeft0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~27 .lut_mask = 16'hBB88;
defparam \ShiftLeft0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N22
cycloneive_lcell_comb \ShiftLeft0~29 (
// Equation(s):
// \ShiftLeft0~29_combout  = (!\Mux92~2_combout  & ((\Mux93~2_combout  & (\ShiftLeft0~110_combout )) # (!\Mux93~2_combout  & ((\ShiftLeft0~28_combout )))))

	.dataa(Mux92),
	.datab(\ShiftLeft0~110_combout ),
	.datac(\ShiftLeft0~28_combout ),
	.datad(Mux931),
	.cin(gnd),
	.combout(\ShiftLeft0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~29 .lut_mask = 16'h4450;
defparam \ShiftLeft0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N0
cycloneive_lcell_comb \ShiftRight0~96 (
// Equation(s):
// \ShiftRight0~96_combout  = (\Mux93~2_combout  & ((\ShiftRight0~33_combout ) # ((\ShiftRight0~34_combout )))) # (!\Mux93~2_combout  & (((\ShiftRight0~55_combout ))))

	.dataa(\ShiftRight0~33_combout ),
	.datab(\ShiftRight0~55_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~34_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~96 .lut_mask = 16'hFCAC;
defparam \ShiftRight0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N10
cycloneive_lcell_comb \portOut~15 (
// Equation(s):
// \portOut~15_combout  = (\Mux24~1_combout  & \Mux88~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux24),
	.datad(Mux88),
	.cin(gnd),
	.combout(\portOut~15_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~15 .lut_mask = 16'hF000;
defparam \portOut~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N6
cycloneive_lcell_comb \aluif.portOut[9]~84 (
// Equation(s):
// \aluif.portOut[9]~84_combout  = (\aluif.portOut[15]~83_combout  & ((\portOut~20_combout ) # ((!\aluif.portOut[15]~82_combout )))) # (!\aluif.portOut[15]~83_combout  & (((\ShiftRight0~105_combout  & \aluif.portOut[15]~82_combout ))))

	.dataa(\aluif.portOut[15]~83_combout ),
	.datab(\portOut~20_combout ),
	.datac(\ShiftRight0~105_combout ),
	.datad(\aluif.portOut[15]~82_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[9]~84_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[9]~84 .lut_mask = 16'hD8AA;
defparam \aluif.portOut[9]~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N10
cycloneive_lcell_comb \portOut~25 (
// Equation(s):
// \portOut~25_combout  = (\Mux23~1_combout  & \Mux87~3_combout )

	.dataa(Mux23),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux87),
	.cin(gnd),
	.combout(\portOut~25_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~25 .lut_mask = 16'hAA00;
defparam \portOut~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y26_N6
cycloneive_lcell_comb \portOut~28 (
// Equation(s):
// \portOut~28_combout  = (\Mux84~3_combout  & \Mux20~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux84),
	.datad(Mux20),
	.cin(gnd),
	.combout(\portOut~28_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~28 .lut_mask = 16'hF000;
defparam \portOut~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N0
cycloneive_lcell_comb \ShiftLeft0~52 (
// Equation(s):
// \ShiftLeft0~52_combout  = (\Mux92~2_combout  & (\ShiftLeft0~21_combout  & (!\Mux93~2_combout ))) # (!\Mux92~2_combout  & (((\ShiftLeft0~51_combout ))))

	.dataa(Mux92),
	.datab(\ShiftLeft0~21_combout ),
	.datac(Mux931),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~52 .lut_mask = 16'h5D08;
defparam \ShiftLeft0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N18
cycloneive_lcell_comb \portOut~31 (
// Equation(s):
// \portOut~31_combout  = (\Mux21~1_combout  & \Mux85~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux21),
	.datad(Mux85),
	.cin(gnd),
	.combout(\portOut~31_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~31 .lut_mask = 16'hF000;
defparam \portOut~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N12
cycloneive_lcell_comb \aluif.portOut[10]~105 (
// Equation(s):
// \aluif.portOut[10]~105_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[15]~26_combout  & \ShiftLeft0~52_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~31_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\portOut~31_combout ),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\ShiftLeft0~52_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[10]~105_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[10]~105 .lut_mask = 16'hE545;
defparam \aluif.portOut[10]~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N26
cycloneive_lcell_comb \portOut~34 (
// Equation(s):
// \portOut~34_combout  = (\Mux18~1_combout  & \Mux82~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux18),
	.datad(Mux82),
	.cin(gnd),
	.combout(\portOut~34_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~34 .lut_mask = 16'hF000;
defparam \portOut~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N10
cycloneive_lcell_comb \ShiftLeft0~61 (
// Equation(s):
// \ShiftLeft0~61_combout  = (\Mux93~2_combout  & ((\ShiftLeft0~42_combout ))) # (!\Mux93~2_combout  & (\ShiftLeft0~60_combout ))

	.dataa(Mux931),
	.datab(gnd),
	.datac(\ShiftLeft0~60_combout ),
	.datad(\ShiftLeft0~42_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~61 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N8
cycloneive_lcell_comb \portOut~37 (
// Equation(s):
// \portOut~37_combout  = (\Mux83~3_combout  & ((\Mux19~1_combout ) # (\Mux19~0_combout )))

	.dataa(Mux191),
	.datab(gnd),
	.datac(Mux83),
	.datad(Mux19),
	.cin(gnd),
	.combout(\portOut~37_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~37 .lut_mask = 16'hF0A0;
defparam \portOut~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N2
cycloneive_lcell_comb \ShiftRight0~111 (
// Equation(s):
// \ShiftRight0~111_combout  = (!\Mux92~2_combout  & (!\ShiftLeft0~5_combout  & \ShiftRight0~43_combout ))

	.dataa(gnd),
	.datab(Mux92),
	.datac(\ShiftLeft0~5_combout ),
	.datad(\ShiftRight0~43_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~111_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~111 .lut_mask = 16'h0300;
defparam \ShiftRight0~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N10
cycloneive_lcell_comb \aluif.portOut[14]~127 (
// Equation(s):
// \aluif.portOut[14]~127_combout  = (\aluif.portOut[15]~82_combout  & ((\aluif.portOut[15]~83_combout  & (\portOut~41_combout )) # (!\aluif.portOut[15]~83_combout  & ((\ShiftRight0~111_combout ))))) # (!\aluif.portOut[15]~82_combout  & 
// (((\aluif.portOut[15]~83_combout ))))

	.dataa(\portOut~41_combout ),
	.datab(\aluif.portOut[15]~82_combout ),
	.datac(\aluif.portOut[15]~83_combout ),
	.datad(\ShiftRight0~111_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[14]~127_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[14]~127 .lut_mask = 16'hBCB0;
defparam \aluif.portOut[14]~127 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N22
cycloneive_lcell_comb \portOut~42 (
// Equation(s):
// \portOut~42_combout  = \Mux81~3_combout  $ (\Mux17~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux81),
	.datad(Mux17),
	.cin(gnd),
	.combout(\portOut~42_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~42 .lut_mask = 16'h0FF0;
defparam \portOut~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N28
cycloneive_lcell_comb \ShiftLeft0~78 (
// Equation(s):
// \ShiftLeft0~78_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout ) # ((\Mux11~1_combout )))) # (!\Mux94~1_combout  & (!\Mux95~1_combout  & ((\Mux9~1_combout ))))

	.dataa(Mux94),
	.datab(Mux95),
	.datac(Mux11),
	.datad(Mux9),
	.cin(gnd),
	.combout(\ShiftLeft0~78_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~78 .lut_mask = 16'hB9A8;
defparam \ShiftLeft0~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N10
cycloneive_lcell_comb \aluif.portOut[29]~157 (
// Equation(s):
// \aluif.portOut[29]~157_combout  = (\aluif.portOut[2]~35_combout  & (((!\ShiftRight0~61_combout )))) # (!\aluif.portOut[2]~35_combout  & ((\ShiftRight0~61_combout  & (\ShiftLeft0~91_combout )) # (!\ShiftRight0~61_combout  & ((\ShiftLeft0~90_combout )))))

	.dataa(\aluif.portOut[2]~35_combout ),
	.datab(\ShiftLeft0~91_combout ),
	.datac(\ShiftLeft0~90_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[29]~157_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~157 .lut_mask = 16'h44FA;
defparam \aluif.portOut[29]~157 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N20
cycloneive_lcell_comb \ShiftLeft0~95 (
// Equation(s):
// \ShiftLeft0~95_combout  = (\Mux95~1_combout  & ((\Mux4~1_combout ))) # (!\Mux95~1_combout  & (\Mux3~1_combout ))

	.dataa(gnd),
	.datab(Mux95),
	.datac(Mux3),
	.datad(Mux4),
	.cin(gnd),
	.combout(\ShiftLeft0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~95 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N26
cycloneive_lcell_comb \aluif.portOut[28]~173 (
// Equation(s):
// \aluif.portOut[28]~173_combout  = (\aluif.portOut[2]~35_combout  & (((!\ShiftRight0~61_combout )))) # (!\aluif.portOut[2]~35_combout  & ((\ShiftRight0~61_combout  & (\ShiftLeft0~95_combout )) # (!\ShiftRight0~61_combout  & ((\ShiftLeft0~94_combout )))))

	.dataa(\aluif.portOut[2]~35_combout ),
	.datab(\ShiftLeft0~95_combout ),
	.datac(\ShiftLeft0~94_combout ),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~173_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~173 .lut_mask = 16'h44FA;
defparam \aluif.portOut[28]~173 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N6
cycloneive_lcell_comb \aluif.portOut[28]~175 (
// Equation(s):
// \aluif.portOut[28]~175_combout  = (\aluif.portOut[1]~13_combout  & ((\aluif.portOut[2]~34_combout  & ((\ShiftLeft0~62_combout ))) # (!\aluif.portOut[2]~34_combout  & (\aluif.portOut[28]~174_combout )))) # (!\aluif.portOut[1]~13_combout  & 
// (((\aluif.portOut[2]~34_combout ))))

	.dataa(\aluif.portOut[28]~174_combout ),
	.datab(\aluif.portOut[1]~13_combout ),
	.datac(\ShiftLeft0~62_combout ),
	.datad(\aluif.portOut[2]~34_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~175_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~175 .lut_mask = 16'hF388;
defparam \aluif.portOut[28]~175 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N18
cycloneive_lcell_comb \portOut~55 (
// Equation(s):
// \portOut~55_combout  = \Mux64~0_combout  $ (\Mux0~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux64),
	.datad(Mux0),
	.cin(gnd),
	.combout(\portOut~55_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~55 .lut_mask = 16'h0FF0;
defparam \portOut~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N4
cycloneive_lcell_comb \portOut~56 (
// Equation(s):
// \portOut~56_combout  = (\Mux0~1_combout  & \Mux64~0_combout )

	.dataa(gnd),
	.datab(Mux0),
	.datac(Mux64),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~56_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~56 .lut_mask = 16'hC0C0;
defparam \portOut~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N14
cycloneive_lcell_comb \aluif.neg_flag~13 (
// Equation(s):
// \aluif.neg_flag~13_combout  = (\aluif.portOut[15]~83_combout  & (((\portOut~56_combout ) # (!\aluif.portOut[15]~82_combout )))) # (!\aluif.portOut[15]~83_combout  & (\ShiftLeft0~67_combout  & ((\aluif.portOut[15]~82_combout ))))

	.dataa(\ShiftLeft0~67_combout ),
	.datab(\aluif.portOut[15]~83_combout ),
	.datac(\portOut~56_combout ),
	.datad(\aluif.portOut[15]~82_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~13_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~13 .lut_mask = 16'hE2CC;
defparam \aluif.neg_flag~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N28
cycloneive_lcell_comb \aluif.portOut[30]~184 (
// Equation(s):
// \aluif.portOut[30]~184_combout  = (\aluif.portOut[30]~181_combout  & (((\ShiftLeft0~5_combout )))) # (!\aluif.portOut[30]~181_combout  & ((\ShiftLeft0~5_combout  & (\ShiftLeft0~95_combout )) # (!\ShiftLeft0~5_combout  & ((\Mux1~1_combout )))))

	.dataa(\aluif.portOut[30]~181_combout ),
	.datab(\ShiftLeft0~95_combout ),
	.datac(\ShiftLeft0~5_combout ),
	.datad(Mux1),
	.cin(gnd),
	.combout(\aluif.portOut[30]~184_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[30]~184 .lut_mask = 16'hE5E0;
defparam \aluif.portOut[30]~184 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N22
cycloneive_lcell_comb \aluif.portOut[30]~185 (
// Equation(s):
// \aluif.portOut[30]~185_combout  = (\aluif.portOut[30]~181_combout  & ((\aluif.portOut[30]~184_combout  & (\ShiftLeft0~104_combout )) # (!\aluif.portOut[30]~184_combout  & ((\Mux2~1_combout ))))) # (!\aluif.portOut[30]~181_combout  & 
// (((\aluif.portOut[30]~184_combout ))))

	.dataa(\ShiftLeft0~104_combout ),
	.datab(\aluif.portOut[30]~181_combout ),
	.datac(Mux2),
	.datad(\aluif.portOut[30]~184_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[30]~185_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[30]~185 .lut_mask = 16'hBBC0;
defparam \aluif.portOut[30]~185 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N10
cycloneive_lcell_comb \portOut~58 (
// Equation(s):
// \portOut~58_combout  = (\Mux65~0_combout  & \Mux1~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux65),
	.datad(Mux1),
	.cin(gnd),
	.combout(\portOut~58_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~58 .lut_mask = 16'hF000;
defparam \portOut~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N10
cycloneive_lcell_comb \aluif.portOut[20]~192 (
// Equation(s):
// \aluif.portOut[20]~192_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & (\ShiftRight0~98_combout )) # (!\prif.ALUOP_ex [2] & ((\portOut~61_combout ))))) # (!\aluif.portOut[15]~26_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\ShiftRight0~98_combout ),
	.datab(\aluif.portOut[15]~26_combout ),
	.datac(prifALUOP_ex_2),
	.datad(\portOut~61_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[20]~192_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[20]~192 .lut_mask = 16'h8F83;
defparam \aluif.portOut[20]~192 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N30
cycloneive_lcell_comb \ShiftLeft0~108 (
// Equation(s):
// \ShiftLeft0~108_combout  = (\Mux93~2_combout  & (\ShiftLeft0~70_combout )) # (!\Mux93~2_combout  & (((\ShiftLeft0~80_combout ) # (\ShiftLeft0~81_combout ))))

	.dataa(\ShiftLeft0~70_combout ),
	.datab(Mux931),
	.datac(\ShiftLeft0~80_combout ),
	.datad(\ShiftLeft0~81_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~108_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~108 .lut_mask = 16'hBBB8;
defparam \ShiftLeft0~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N18
cycloneive_lcell_comb \aluif.portOut[18]~216 (
// Equation(s):
// \aluif.portOut[18]~216_combout  = (\ShiftLeft0~108_combout  & (((!\aluif.portOut[15]~83_combout )))) # (!\ShiftLeft0~108_combout  & (\aluif.portOut[15]~82_combout  & ((\ShiftLeft0~109_combout ) # (\aluif.portOut[15]~83_combout ))))

	.dataa(\ShiftLeft0~109_combout ),
	.datab(\aluif.portOut[15]~82_combout ),
	.datac(\aluif.portOut[15]~83_combout ),
	.datad(\ShiftLeft0~108_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[18]~216_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[18]~216 .lut_mask = 16'h0FC8;
defparam \aluif.portOut[18]~216 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N12
cycloneive_lcell_comb \aluif.portOut[18]~217 (
// Equation(s):
// \aluif.portOut[18]~217_combout  = (\aluif.portOut[15]~83_combout  & (((\Mux77~0_combout  & \Mux13~1_combout )) # (!\aluif.portOut[18]~216_combout ))) # (!\aluif.portOut[15]~83_combout  & (((\aluif.portOut[18]~216_combout ))))

	.dataa(\aluif.portOut[15]~83_combout ),
	.datab(Mux77),
	.datac(Mux13),
	.datad(\aluif.portOut[18]~216_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[18]~217_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[18]~217 .lut_mask = 16'hD5AA;
defparam \aluif.portOut[18]~217 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N12
cycloneive_lcell_comb \aluif.portOut[27]~242 (
// Equation(s):
// \aluif.portOut[27]~242_combout  = (\aluif.portOut[5]~52_combout  & ((\aluif.portOut[5]~51_combout ) # ((\ShiftLeft0~74_combout )))) # (!\aluif.portOut[5]~52_combout  & (!\aluif.portOut[5]~51_combout  & (\ShiftLeft0~102_combout )))

	.dataa(\aluif.portOut[5]~52_combout ),
	.datab(\aluif.portOut[5]~51_combout ),
	.datac(\ShiftLeft0~102_combout ),
	.datad(\ShiftLeft0~74_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[27]~242_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[27]~242 .lut_mask = 16'hBA98;
defparam \aluif.portOut[27]~242 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N30
cycloneive_lcell_comb \aluif.portOut[27]~243 (
// Equation(s):
// \aluif.portOut[27]~243_combout  = (\aluif.portOut[27]~242_combout  & ((\ShiftLeft0~48_combout ) # ((!\aluif.portOut[5]~51_combout )))) # (!\aluif.portOut[27]~242_combout  & (((\aluif.portOut[5]~51_combout  & \ShiftLeft0~107_combout ))))

	.dataa(\aluif.portOut[27]~242_combout ),
	.datab(\ShiftLeft0~48_combout ),
	.datac(\aluif.portOut[5]~51_combout ),
	.datad(\ShiftLeft0~107_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[27]~243_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[27]~243 .lut_mask = 16'hDA8A;
defparam \aluif.portOut[27]~243 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N30
cycloneive_lcell_comb \aluif.neg_flag~23 (
// Equation(s):
// \aluif.neg_flag~23_combout  = ((!\portOut~55_combout  & (!\prif.ALUOP_ex [1] & !\prif.ALUOP_ex [2]))) # (!\prif.ALUOP_ex [0])

	.dataa(prifALUOP_ex_0),
	.datab(\portOut~55_combout ),
	.datac(prifALUOP_ex_1),
	.datad(prifALUOP_ex_2),
	.cin(gnd),
	.combout(\aluif.neg_flag~23_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~23 .lut_mask = 16'h5557;
defparam \aluif.neg_flag~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N22
cycloneive_lcell_comb \aluif.portOut[1]~15 (
// Equation(s):
// aluifportOut_1 = (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [0] & (\aluif.portOut[1]~10_combout )) # (!\prif.ALUOP_ex [0] & ((\aluif.portOut[1]~14_combout )))))

	.dataa(prifALUOP_ex_3),
	.datab(\aluif.portOut[1]~10_combout ),
	.datac(prifALUOP_ex_0),
	.datad(\aluif.portOut[1]~14_combout ),
	.cin(gnd),
	.combout(aluifportOut_1),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[1]~15 .lut_mask = 16'h8A80;
defparam \aluif.portOut[1]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N22
cycloneive_lcell_comb \aluif.portOut[0]~24 (
// Equation(s):
// aluifportOut_0 = (\aluif.portOut[0]~22_combout ) # ((!\prif.ALUOP_ex [1] & (!\prif.ALUOP_ex [3] & \aluif.portOut[0]~23_combout )))

	.dataa(prifALUOP_ex_1),
	.datab(prifALUOP_ex_3),
	.datac(\aluif.portOut[0]~22_combout ),
	.datad(\aluif.portOut[0]~23_combout ),
	.cin(gnd),
	.combout(aluifportOut_0),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[0]~24 .lut_mask = 16'hF1F0;
defparam \aluif.portOut[0]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N8
cycloneive_lcell_comb \aluif.portOut[3]~30 (
// Equation(s):
// aluifportOut_3 = (\portOut~4_combout  & (\aluif.portOut[5]~25_combout  & ((\aluif.portOut[3]~28_combout )))) # (!\portOut~4_combout  & ((\aluif.portOut[2]~29_combout ) # ((\aluif.portOut[5]~25_combout  & \aluif.portOut[3]~28_combout ))))

	.dataa(\portOut~4_combout ),
	.datab(\aluif.portOut[5]~25_combout ),
	.datac(\aluif.portOut[2]~29_combout ),
	.datad(\aluif.portOut[3]~28_combout ),
	.cin(gnd),
	.combout(aluifportOut_3),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[3]~30 .lut_mask = 16'hDC50;
defparam \aluif.portOut[3]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N8
cycloneive_lcell_comb \aluif.portOut[5]~31 (
// Equation(s):
// aluifportOut_5 = (!\prif.ALUOP_ex [0] & \prif.ALUOP_ex [3])

	.dataa(gnd),
	.datab(prifALUOP_ex_0),
	.datac(prifALUOP_ex_3),
	.datad(gnd),
	.cin(gnd),
	.combout(aluifportOut_5),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~31 .lut_mask = 16'h3030;
defparam \aluif.portOut[5]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N14
cycloneive_lcell_comb \aluif.portOut[2]~33 (
// Equation(s):
// aluifportOut_2 = (aluifportOut_5 & (!\aluif.portOut[2]~32_combout  & ((!\ShiftLeft0~15_combout ) # (!\aluif.portOut[1]~13_combout ))))

	.dataa(aluifportOut_5),
	.datab(\aluif.portOut[1]~13_combout ),
	.datac(\aluif.portOut[2]~32_combout ),
	.datad(\ShiftLeft0~15_combout ),
	.cin(gnd),
	.combout(aluifportOut_2),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~33 .lut_mask = 16'h020A;
defparam \aluif.portOut[2]~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N6
cycloneive_lcell_comb \aluif.portOut[3]~39 (
// Equation(s):
// aluifportOut_31 = (\aluif.portOut[1]~13_combout  & (((\aluif.portOut[3]~38_combout )))) # (!\aluif.portOut[1]~13_combout  & ((\aluif.portOut[3]~38_combout  & (\Add1~6_combout )) # (!\aluif.portOut[3]~38_combout  & ((\portOut~4_combout )))))

	.dataa(\aluif.portOut[1]~13_combout ),
	.datab(\Add1~6_combout ),
	.datac(\portOut~4_combout ),
	.datad(\aluif.portOut[3]~38_combout ),
	.cin(gnd),
	.combout(aluifportOut_31),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[3]~39 .lut_mask = 16'hEE50;
defparam \aluif.portOut[3]~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N28
cycloneive_lcell_comb \aluif.portOut[3]~40 (
// Equation(s):
// aluifportOut_32 = (aluifportOut_3) # ((aluifportOut_2 & aluifportOut_31))

	.dataa(gnd),
	.datab(aluifportOut_2),
	.datac(aluifportOut_3),
	.datad(aluifportOut_31),
	.cin(gnd),
	.combout(aluifportOut_32),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[3]~40 .lut_mask = 16'hFCF0;
defparam \aluif.portOut[3]~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N12
cycloneive_lcell_comb \aluif.portOut[2]~48 (
// Equation(s):
// aluifportOut_21 = (\aluif.portOut[2]~43_combout ) # ((\aluif.portOut[2]~47_combout  & aluifportOut_2))

	.dataa(gnd),
	.datab(\aluif.portOut[2]~47_combout ),
	.datac(aluifportOut_2),
	.datad(\aluif.portOut[2]~43_combout ),
	.cin(gnd),
	.combout(aluifportOut_21),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~48 .lut_mask = 16'hFFC0;
defparam \aluif.portOut[2]~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N4
cycloneive_lcell_comb \aluif.portOut[5]~57 (
// Equation(s):
// aluifportOut_51 = (\aluif.portOut[5]~56_combout  & (((\prif.ALUOP_ex [1]) # (!\portOut~10_combout )))) # (!\aluif.portOut[5]~56_combout  & (\Add1~10_combout  & ((!\prif.ALUOP_ex [1]))))

	.dataa(\Add1~10_combout ),
	.datab(\portOut~10_combout ),
	.datac(\aluif.portOut[5]~56_combout ),
	.datad(prifALUOP_ex_1),
	.cin(gnd),
	.combout(aluifportOut_51),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~57 .lut_mask = 16'hF03A;
defparam \aluif.portOut[5]~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N16
cycloneive_lcell_comb \aluif.portOut[5]~58 (
// Equation(s):
// aluifportOut_52 = (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [0] & ((\aluif.portOut[5]~50_combout ))) # (!\prif.ALUOP_ex [0] & (aluifportOut_51))))

	.dataa(prifALUOP_ex_3),
	.datab(aluifportOut_51),
	.datac(prifALUOP_ex_0),
	.datad(\aluif.portOut[5]~50_combout ),
	.cin(gnd),
	.combout(aluifportOut_52),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~58 .lut_mask = 16'hA808;
defparam \aluif.portOut[5]~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N0
cycloneive_lcell_comb \aluif.portOut[4]~65 (
// Equation(s):
// aluifportOut_4 = (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [0] & (\aluif.portOut[4]~60_combout )) # (!\prif.ALUOP_ex [0] & ((\aluif.portOut[4]~64_combout )))))

	.dataa(prifALUOP_ex_0),
	.datab(prifALUOP_ex_3),
	.datac(\aluif.portOut[4]~60_combout ),
	.datad(\aluif.portOut[4]~64_combout ),
	.cin(gnd),
	.combout(aluifportOut_4),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[4]~65 .lut_mask = 16'hC480;
defparam \aluif.portOut[4]~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N22
cycloneive_lcell_comb \aluif.portOut[7]~72 (
// Equation(s):
// aluifportOut_7 = (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [0] & ((\aluif.portOut[7]~67_combout ))) # (!\prif.ALUOP_ex [0] & (\aluif.portOut[7]~71_combout ))))

	.dataa(prifALUOP_ex_0),
	.datab(prifALUOP_ex_3),
	.datac(\aluif.portOut[7]~71_combout ),
	.datad(\aluif.portOut[7]~67_combout ),
	.cin(gnd),
	.combout(aluifportOut_7),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[7]~72 .lut_mask = 16'hC840;
defparam \aluif.portOut[7]~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N26
cycloneive_lcell_comb \aluif.portOut[6]~79 (
// Equation(s):
// aluifportOut_6 = (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [0] & (\aluif.portOut[6]~74_combout )) # (!\prif.ALUOP_ex [0] & ((\aluif.portOut[6]~78_combout )))))

	.dataa(prifALUOP_ex_0),
	.datab(prifALUOP_ex_3),
	.datac(\aluif.portOut[6]~74_combout ),
	.datad(\aluif.portOut[6]~78_combout ),
	.cin(gnd),
	.combout(aluifportOut_6),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[6]~79 .lut_mask = 16'hC480;
defparam \aluif.portOut[6]~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N24
cycloneive_lcell_comb \aluif.portOut[9]~90 (
// Equation(s):
// aluifportOut_9 = (\aluif.portOut[15]~80_combout  & ((\aluif.portOut[9]~89_combout  & ((!\portOut~20_combout ))) # (!\aluif.portOut[9]~89_combout  & (\Add1~18_combout )))) # (!\aluif.portOut[15]~80_combout  & (((\aluif.portOut[9]~89_combout ))))

	.dataa(\Add1~18_combout ),
	.datab(\aluif.portOut[15]~80_combout ),
	.datac(\aluif.portOut[9]~89_combout ),
	.datad(\portOut~20_combout ),
	.cin(gnd),
	.combout(aluifportOut_9),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[9]~90 .lut_mask = 16'h38F8;
defparam \aluif.portOut[9]~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N18
cycloneive_lcell_comb \aluif.portOut[8]~96 (
// Equation(s):
// aluifportOut_8 = (\aluif.portOut[8]~95_combout  & (((!\aluif.portOut[15]~86_combout )) # (!\portOut~23_combout ))) # (!\aluif.portOut[8]~95_combout  & (((\aluif.portOut[8]~92_combout  & \aluif.portOut[15]~86_combout ))))

	.dataa(\portOut~23_combout ),
	.datab(\aluif.portOut[8]~95_combout ),
	.datac(\aluif.portOut[8]~92_combout ),
	.datad(\aluif.portOut[15]~86_combout ),
	.cin(gnd),
	.combout(aluifportOut_8),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[8]~96 .lut_mask = 16'h74CC;
defparam \aluif.portOut[8]~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N6
cycloneive_lcell_comb \aluif.portOut[11]~102 (
// Equation(s):
// aluifportOut_11 = (\aluif.portOut[11]~101_combout  & (((!\aluif.portOut[15]~80_combout )) # (!\portOut~26_combout ))) # (!\aluif.portOut[11]~101_combout  & (((\aluif.portOut[15]~80_combout  & \Add1~22_combout ))))

	.dataa(\portOut~26_combout ),
	.datab(\aluif.portOut[11]~101_combout ),
	.datac(\aluif.portOut[15]~80_combout ),
	.datad(\Add1~22_combout ),
	.cin(gnd),
	.combout(aluifportOut_11),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[11]~102 .lut_mask = 16'h7C4C;
defparam \aluif.portOut[11]~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N2
cycloneive_lcell_comb \aluif.portOut[10]~108 (
// Equation(s):
// aluifportOut_10 = (\aluif.portOut[10]~107_combout  & (((!\aluif.portOut[15]~86_combout )) # (!\portOut~29_combout ))) # (!\aluif.portOut[10]~107_combout  & (((\aluif.portOut[15]~86_combout  & \aluif.portOut[10]~104_combout ))))

	.dataa(\portOut~29_combout ),
	.datab(\aluif.portOut[10]~107_combout ),
	.datac(\aluif.portOut[15]~86_combout ),
	.datad(\aluif.portOut[10]~104_combout ),
	.cin(gnd),
	.combout(aluifportOut_10),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[10]~108 .lut_mask = 16'h7C4C;
defparam \aluif.portOut[10]~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N22
cycloneive_lcell_comb \aluif.portOut[13]~114 (
// Equation(s):
// aluifportOut_13 = (\aluif.portOut[15]~86_combout  & ((\aluif.portOut[13]~113_combout  & ((!\portOut~32_combout ))) # (!\aluif.portOut[13]~113_combout  & (\aluif.portOut[13]~110_combout )))) # (!\aluif.portOut[15]~86_combout  & 
// (((\aluif.portOut[13]~113_combout ))))

	.dataa(\aluif.portOut[13]~110_combout ),
	.datab(\portOut~32_combout ),
	.datac(\aluif.portOut[15]~86_combout ),
	.datad(\aluif.portOut[13]~113_combout ),
	.cin(gnd),
	.combout(aluifportOut_13),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[13]~114 .lut_mask = 16'h3FA0;
defparam \aluif.portOut[13]~114 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N4
cycloneive_lcell_comb \aluif.portOut[12]~120 (
// Equation(s):
// aluifportOut_12 = (\aluif.portOut[15]~80_combout  & ((\aluif.portOut[12]~119_combout  & ((!\portOut~35_combout ))) # (!\aluif.portOut[12]~119_combout  & (\Add1~24_combout )))) # (!\aluif.portOut[15]~80_combout  & (((\aluif.portOut[12]~119_combout ))))

	.dataa(\Add1~24_combout ),
	.datab(\portOut~35_combout ),
	.datac(\aluif.portOut[15]~80_combout ),
	.datad(\aluif.portOut[12]~119_combout ),
	.cin(gnd),
	.combout(aluifportOut_12),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[12]~120 .lut_mask = 16'h3FA0;
defparam \aluif.portOut[12]~120 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N26
cycloneive_lcell_comb \aluif.portOut[15]~126 (
// Equation(s):
// aluifportOut_15 = (\aluif.portOut[15]~86_combout  & ((\aluif.portOut[15]~125_combout  & (!\portOut~38_combout )) # (!\aluif.portOut[15]~125_combout  & ((\aluif.portOut[15]~122_combout ))))) # (!\aluif.portOut[15]~86_combout  & 
// (((\aluif.portOut[15]~125_combout ))))

	.dataa(\portOut~38_combout ),
	.datab(\aluif.portOut[15]~86_combout ),
	.datac(\aluif.portOut[15]~125_combout ),
	.datad(\aluif.portOut[15]~122_combout ),
	.cin(gnd),
	.combout(aluifportOut_15),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~126 .lut_mask = 16'h7C70;
defparam \aluif.portOut[15]~126 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N0
cycloneive_lcell_comb \aluif.portOut[14]~132 (
// Equation(s):
// aluifportOut_14 = (\aluif.portOut[15]~80_combout  & ((\aluif.portOut[14]~131_combout  & ((!\portOut~41_combout ))) # (!\aluif.portOut[14]~131_combout  & (\Add1~28_combout )))) # (!\aluif.portOut[15]~80_combout  & (((\aluif.portOut[14]~131_combout ))))

	.dataa(\Add1~28_combout ),
	.datab(\aluif.portOut[15]~80_combout ),
	.datac(\portOut~41_combout ),
	.datad(\aluif.portOut[14]~131_combout ),
	.cin(gnd),
	.combout(aluifportOut_14),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[14]~132 .lut_mask = 16'h3F88;
defparam \aluif.portOut[14]~132 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N30
cycloneive_lcell_comb \aluif.portOut[23]~140 (
// Equation(s):
// aluifportOut_23 = (\aluif.portOut[23]~135_combout  & ((\aluif.portOut[23]~139_combout  & ((\portOut~46_combout ))) # (!\aluif.portOut[23]~139_combout  & (\aluif.portOut[23]~134_combout )))) # (!\aluif.portOut[23]~135_combout  & 
// (((\aluif.portOut[23]~139_combout ))))

	.dataa(\aluif.portOut[23]~134_combout ),
	.datab(\portOut~46_combout ),
	.datac(\aluif.portOut[23]~135_combout ),
	.datad(\aluif.portOut[23]~139_combout ),
	.cin(gnd),
	.combout(aluifportOut_23),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[23]~140 .lut_mask = 16'hCFA0;
defparam \aluif.portOut[23]~140 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N28
cycloneive_lcell_comb \aluif.portOut[22]~147 (
// Equation(s):
// aluifportOut_22 = (\aluif.portOut[22]~145_combout  & ((\Add0~44_combout ) # ((\aluif.portOut[22]~261_combout )))) # (!\aluif.portOut[22]~145_combout  & (((\Add1~44_combout  & \aluif.portOut[22]~261_combout ))))

	.dataa(\aluif.portOut[22]~145_combout ),
	.datab(\Add0~44_combout ),
	.datac(\Add1~44_combout ),
	.datad(\aluif.portOut[22]~261_combout ),
	.cin(gnd),
	.combout(aluifportOut_22),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~147 .lut_mask = 16'hFA88;
defparam \aluif.portOut[22]~147 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N14
cycloneive_lcell_comb \aluif.portOut[21]~153 (
// Equation(s):
// aluifportOut_211 = (\aluif.portOut[23]~135_combout  & ((\aluif.portOut[21]~152_combout  & (\portOut~51_combout )) # (!\aluif.portOut[21]~152_combout  & ((\aluif.portOut[21]~149_combout ))))) # (!\aluif.portOut[23]~135_combout  & 
// (((\aluif.portOut[21]~152_combout ))))

	.dataa(\portOut~51_combout ),
	.datab(\aluif.portOut[23]~135_combout ),
	.datac(\aluif.portOut[21]~149_combout ),
	.datad(\aluif.portOut[21]~152_combout ),
	.cin(gnd),
	.combout(aluifportOut_211),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[21]~153 .lut_mask = 16'hBBC0;
defparam \aluif.portOut[21]~153 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N2
cycloneive_lcell_comb \aluif.portOut[29]~166 (
// Equation(s):
// aluifportOut_29 = (\aluif.portOut[29]~165_combout ) # ((\aluif.portOut[29]~161_combout ) # ((\aluif.portOut[28]~154_combout  & \aluif.portOut[29]~162_combout )))

	.dataa(\aluif.portOut[28]~154_combout ),
	.datab(\aluif.portOut[29]~165_combout ),
	.datac(\aluif.portOut[29]~162_combout ),
	.datad(\aluif.portOut[29]~161_combout ),
	.cin(gnd),
	.combout(aluifportOut_29),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~166 .lut_mask = 16'hFFEC;
defparam \aluif.portOut[29]~166 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N12
cycloneive_lcell_comb \aluif.portOut[28]~180 (
// Equation(s):
// aluifportOut_28 = (\aluif.portOut[28]~179_combout ) # ((\aluif.portOut[28]~167_combout ) # ((\aluif.portOut[28]~170_combout  & \Add1~56_combout )))

	.dataa(\aluif.portOut[28]~179_combout ),
	.datab(\aluif.portOut[28]~167_combout ),
	.datac(\aluif.portOut[28]~170_combout ),
	.datad(\Add1~56_combout ),
	.cin(gnd),
	.combout(aluifportOut_28),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~180 .lut_mask = 16'hFEEE;
defparam \aluif.portOut[28]~180 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N26
cycloneive_lcell_comb \aluif.neg_flag~19 (
// Equation(s):
// aluifneg_flag = (\aluif.neg_flag~22_combout  & (((\Add1~62_combout ) # (\aluif.neg_flag~17_combout )))) # (!\aluif.neg_flag~22_combout  & (\Add0~62_combout  & ((\aluif.neg_flag~17_combout ))))

	.dataa(\Add0~62_combout ),
	.datab(\Add1~62_combout ),
	.datac(\aluif.neg_flag~22_combout ),
	.datad(\aluif.neg_flag~17_combout ),
	.cin(gnd),
	.combout(aluifneg_flag),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~19 .lut_mask = 16'hFAC0;
defparam \aluif.neg_flag~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N0
cycloneive_lcell_comb \aluif.portOut[30]~189 (
// Equation(s):
// aluifportOut_30 = (\aluif.portOut[23]~135_combout  & ((\aluif.portOut[30]~188_combout  & (\portOut~59_combout )) # (!\aluif.portOut[30]~188_combout  & ((\aluif.portOut[30]~183_combout ))))) # (!\aluif.portOut[23]~135_combout  & 
// (((\aluif.portOut[30]~188_combout ))))

	.dataa(\aluif.portOut[23]~135_combout ),
	.datab(\portOut~59_combout ),
	.datac(\aluif.portOut[30]~183_combout ),
	.datad(\aluif.portOut[30]~188_combout ),
	.cin(gnd),
	.combout(aluifportOut_30),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[30]~189 .lut_mask = 16'hDDA0;
defparam \aluif.portOut[30]~189 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N30
cycloneive_lcell_comb \aluif.portOut[20]~195 (
// Equation(s):
// aluifportOut_20 = (\aluif.portOut[23]~136_combout  & ((\aluif.portOut[20]~194_combout  & (\portOut~62_combout )) # (!\aluif.portOut[20]~194_combout  & ((\Add0~40_combout ))))) # (!\aluif.portOut[23]~136_combout  & (((\aluif.portOut[20]~194_combout ))))

	.dataa(\aluif.portOut[23]~136_combout ),
	.datab(\portOut~62_combout ),
	.datac(\Add0~40_combout ),
	.datad(\aluif.portOut[20]~194_combout ),
	.cin(gnd),
	.combout(aluifportOut_20),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[20]~195 .lut_mask = 16'hDDA0;
defparam \aluif.portOut[20]~195 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N22
cycloneive_lcell_comb \aluif.portOut[17]~201 (
// Equation(s):
// aluifportOut_17 = (\aluif.portOut[23]~136_combout  & ((\aluif.portOut[17]~200_combout  & ((\portOut~65_combout ))) # (!\aluif.portOut[17]~200_combout  & (\Add0~34_combout )))) # (!\aluif.portOut[23]~136_combout  & (((\aluif.portOut[17]~200_combout ))))

	.dataa(\Add0~34_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(\portOut~65_combout ),
	.datad(\aluif.portOut[17]~200_combout ),
	.cin(gnd),
	.combout(aluifportOut_17),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[17]~201 .lut_mask = 16'hF388;
defparam \aluif.portOut[17]~201 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y25_N2
cycloneive_lcell_comb \aluif.portOut[16]~207 (
// Equation(s):
// aluifportOut_16 = (\aluif.portOut[16]~206_combout  & ((\portOut~68_combout ) # ((!\aluif.portOut[23]~135_combout )))) # (!\aluif.portOut[16]~206_combout  & (((\aluif.portOut[23]~135_combout  & \aluif.portOut[16]~203_combout ))))

	.dataa(\aluif.portOut[16]~206_combout ),
	.datab(\portOut~68_combout ),
	.datac(\aluif.portOut[23]~135_combout ),
	.datad(\aluif.portOut[16]~203_combout ),
	.cin(gnd),
	.combout(aluifportOut_16),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[16]~207 .lut_mask = 16'hDA8A;
defparam \aluif.portOut[16]~207 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N10
cycloneive_lcell_comb \aluif.portOut[19]~213 (
// Equation(s):
// aluifportOut_19 = (\aluif.portOut[23]~135_combout  & ((\aluif.portOut[19]~212_combout  & (\portOut~71_combout )) # (!\aluif.portOut[19]~212_combout  & ((\aluif.portOut[19]~209_combout ))))) # (!\aluif.portOut[23]~135_combout  & 
// (((\aluif.portOut[19]~212_combout ))))

	.dataa(\portOut~71_combout ),
	.datab(\aluif.portOut[23]~135_combout ),
	.datac(\aluif.portOut[19]~212_combout ),
	.datad(\aluif.portOut[19]~209_combout ),
	.cin(gnd),
	.combout(aluifportOut_19),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[19]~213 .lut_mask = 16'hBCB0;
defparam \aluif.portOut[19]~213 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N16
cycloneive_lcell_comb \aluif.portOut[18]~221 (
// Equation(s):
// aluifportOut_18 = (\aluif.portOut[23]~136_combout  & ((\aluif.portOut[18]~220_combout  & (\portOut~74_combout )) # (!\aluif.portOut[18]~220_combout  & ((\Add0~36_combout ))))) # (!\aluif.portOut[23]~136_combout  & (((\aluif.portOut[18]~220_combout ))))

	.dataa(\portOut~74_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(\Add0~36_combout ),
	.datad(\aluif.portOut[18]~220_combout ),
	.cin(gnd),
	.combout(aluifportOut_18),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[18]~221 .lut_mask = 16'hBBC0;
defparam \aluif.portOut[18]~221 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N24
cycloneive_lcell_comb \aluif.portOut[25]~234 (
// Equation(s):
// aluifportOut_25 = (\aluif.portOut[25]~233_combout  & (((\Add0~50_combout ) # (\aluif.portOut[25]~224_combout )) # (!\prif.ALUOP_ex [0])))

	.dataa(\aluif.portOut[25]~233_combout ),
	.datab(prifALUOP_ex_0),
	.datac(\Add0~50_combout ),
	.datad(\aluif.portOut[25]~224_combout ),
	.cin(gnd),
	.combout(aluifportOut_25),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~234 .lut_mask = 16'hAAA2;
defparam \aluif.portOut[25]~234 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N16
cycloneive_lcell_comb \aluif.portOut[24]~241 (
// Equation(s):
// aluifportOut_24 = (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [0] & (\aluif.portOut[24]~238_combout )) # (!\prif.ALUOP_ex [0] & ((\aluif.portOut[24]~240_combout )))))

	.dataa(prifALUOP_ex_3),
	.datab(prifALUOP_ex_0),
	.datac(\aluif.portOut[24]~238_combout ),
	.datad(\aluif.portOut[24]~240_combout ),
	.cin(gnd),
	.combout(aluifportOut_24),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[24]~241 .lut_mask = 16'hA280;
defparam \aluif.portOut[24]~241 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N14
cycloneive_lcell_comb \aluif.portOut[27]~249 (
// Equation(s):
// aluifportOut_27 = (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [0] & ((\aluif.portOut[27]~246_combout ))) # (!\prif.ALUOP_ex [0] & (\aluif.portOut[27]~248_combout ))))

	.dataa(prifALUOP_ex_0),
	.datab(\aluif.portOut[27]~248_combout ),
	.datac(prifALUOP_ex_3),
	.datad(\aluif.portOut[27]~246_combout ),
	.cin(gnd),
	.combout(aluifportOut_27),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[27]~249 .lut_mask = 16'hE040;
defparam \aluif.portOut[27]~249 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N14
cycloneive_lcell_comb \aluif.portOut[26]~257 (
// Equation(s):
// aluifportOut_26 = (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [0] & ((\aluif.portOut[26]~254_combout ))) # (!\prif.ALUOP_ex [0] & (\aluif.portOut[26]~256_combout ))))

	.dataa(\aluif.portOut[26]~256_combout ),
	.datab(prifALUOP_ex_0),
	.datac(prifALUOP_ex_3),
	.datad(\aluif.portOut[26]~254_combout ),
	.cin(gnd),
	.combout(aluifportOut_26),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[26]~257 .lut_mask = 16'hE020;
defparam \aluif.portOut[26]~257 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N18
cycloneive_lcell_comb \aluif.portOut[5]~258 (
// Equation(s):
// aluifportOut_53 = (\prif.ALUOP_ex [3] & (\aluif.portOut[5]~50_combout  & \prif.ALUOP_ex [0]))

	.dataa(prifALUOP_ex_3),
	.datab(\aluif.portOut[5]~50_combout ),
	.datac(gnd),
	.datad(prifALUOP_ex_0),
	.cin(gnd),
	.combout(aluifportOut_53),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~258 .lut_mask = 16'h8800;
defparam \aluif.portOut[5]~258 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N14
cycloneive_lcell_comb \aluif.portOut[1]~9 (
// Equation(s):
// \aluif.portOut[1]~9_combout  = (\prif.ALUOP_ex [2] & (\prif.ALUOP_ex [1])) # (!\prif.ALUOP_ex [2] & ((\prif.ALUOP_ex [1] & (\Mux94~1_combout  & \Mux30~1_combout )) # (!\prif.ALUOP_ex [1] & (\Mux94~1_combout  $ (\Mux30~1_combout )))))

	.dataa(prifALUOP_ex_2),
	.datab(prifALUOP_ex_1),
	.datac(Mux94),
	.datad(Mux30),
	.cin(gnd),
	.combout(\aluif.portOut[1]~9_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[1]~9 .lut_mask = 16'hC998;
defparam \aluif.portOut[1]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N20
cycloneive_lcell_comb \ShiftLeft0~9 (
// Equation(s):
// \ShiftLeft0~9_combout  = (\Mux84~3_combout ) # ((\Mux85~3_combout ) # ((\Mux83~3_combout ) # (\Mux86~3_combout )))

	.dataa(Mux84),
	.datab(Mux85),
	.datac(Mux83),
	.datad(Mux86),
	.cin(gnd),
	.combout(\ShiftLeft0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~9 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N24
cycloneive_lcell_comb \ShiftLeft0~11 (
// Equation(s):
// \ShiftLeft0~11_combout  = (\Mux71~0_combout ) # ((\Mux79~0_combout ) # ((\Mux76~0_combout ) # (\Mux78~0_combout )))

	.dataa(Mux71),
	.datab(Mux79),
	.datac(Mux76),
	.datad(Mux78),
	.cin(gnd),
	.combout(\ShiftLeft0~11_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~11 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N14
cycloneive_lcell_comb \ShiftLeft0~10 (
// Equation(s):
// \ShiftLeft0~10_combout  = (\Mux77~0_combout ) # ((\Mux89~4_combout ) # ((\Mux72~0_combout ) # (\Mux68~0_combout )))

	.dataa(Mux77),
	.datab(Mux891),
	.datac(Mux72),
	.datad(Mux68),
	.cin(gnd),
	.combout(\ShiftLeft0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~10 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N28
cycloneive_lcell_comb \ShiftLeft0~13 (
// Equation(s):
// \ShiftLeft0~13_combout  = (\Mux73~0_combout ) # ((\Mux87~3_combout ) # ((\Mux70~0_combout ) # (\Mux88~3_combout )))

	.dataa(Mux73),
	.datab(Mux87),
	.datac(Mux70),
	.datad(Mux88),
	.cin(gnd),
	.combout(\ShiftLeft0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~13 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N26
cycloneive_lcell_comb \ShiftLeft0~14 (
// Equation(s):
// \ShiftLeft0~14_combout  = (\ShiftLeft0~12_combout ) # ((\ShiftLeft0~11_combout ) # ((\ShiftLeft0~10_combout ) # (\ShiftLeft0~13_combout )))

	.dataa(\ShiftLeft0~12_combout ),
	.datab(\ShiftLeft0~11_combout ),
	.datac(\ShiftLeft0~10_combout ),
	.datad(\ShiftLeft0~13_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~14 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N12
cycloneive_lcell_comb \ShiftLeft0~7 (
// Equation(s):
// \ShiftLeft0~7_combout  = (\Mux64~0_combout ) # ((\Mux66~0_combout ) # (\Mux65~0_combout ))

	.dataa(Mux64),
	.datab(gnd),
	.datac(Mux66),
	.datad(Mux65),
	.cin(gnd),
	.combout(\ShiftLeft0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~7 .lut_mask = 16'hFFFA;
defparam \ShiftLeft0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N4
cycloneive_lcell_comb \ShiftLeft0~15 (
// Equation(s):
// \ShiftLeft0~15_combout  = (\ShiftLeft0~8_combout ) # ((\ShiftLeft0~9_combout ) # ((\ShiftLeft0~14_combout ) # (\ShiftLeft0~7_combout )))

	.dataa(\ShiftLeft0~8_combout ),
	.datab(\ShiftLeft0~9_combout ),
	.datac(\ShiftLeft0~14_combout ),
	.datad(\ShiftLeft0~7_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~15 .lut_mask = 16'hFFFE;
defparam \ShiftLeft0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N8
cycloneive_lcell_comb \ShiftLeft0~5 (
// Equation(s):
// \ShiftLeft0~5_combout  = (\Mux93~0_combout ) # ((\Mux94~1_combout ) # ((\Mux89~2_combout  & \Mux61~1_combout )))

	.dataa(Mux93),
	.datab(Mux89),
	.datac(Mux61),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftLeft0~5_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~5 .lut_mask = 16'hFFEA;
defparam \ShiftLeft0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N8
cycloneive_lcell_comb \ShiftLeft0~4 (
// Equation(s):
// \ShiftLeft0~4_combout  = (\Mux95~1_combout  & (\Mux31~1_combout )) # (!\Mux95~1_combout  & ((\Mux30~1_combout )))

	.dataa(gnd),
	.datab(Mux95),
	.datac(Mux31),
	.datad(Mux30),
	.cin(gnd),
	.combout(\ShiftLeft0~4_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~4 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y22_N16
cycloneive_lcell_comb \ShiftLeft0~6 (
// Equation(s):
// \ShiftLeft0~6_combout  = (!\Mux92~2_combout  & (!\ShiftLeft0~5_combout  & \ShiftLeft0~4_combout ))

	.dataa(gnd),
	.datab(Mux92),
	.datac(\ShiftLeft0~5_combout ),
	.datad(\ShiftLeft0~4_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~6 .lut_mask = 16'h0300;
defparam \ShiftLeft0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N8
cycloneive_lcell_comb \aluif.portOut[1]~8 (
// Equation(s):
// \aluif.portOut[1]~8_combout  = (!\Mux91~2_combout  & (!\ShiftLeft0~15_combout  & \ShiftLeft0~6_combout ))

	.dataa(Mux91),
	.datab(\ShiftLeft0~15_combout ),
	.datac(\ShiftLeft0~6_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\aluif.portOut[1]~8_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[1]~8 .lut_mask = 16'h1010;
defparam \aluif.portOut[1]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N2
cycloneive_lcell_comb \Add0~2 (
// Equation(s):
// \Add0~2_combout  = (\Mux94~1_combout  & ((\Mux30~1_combout  & (\Add0~1  & VCC)) # (!\Mux30~1_combout  & (!\Add0~1 )))) # (!\Mux94~1_combout  & ((\Mux30~1_combout  & (!\Add0~1 )) # (!\Mux30~1_combout  & ((\Add0~1 ) # (GND)))))
// \Add0~3  = CARRY((\Mux94~1_combout  & (!\Mux30~1_combout  & !\Add0~1 )) # (!\Mux94~1_combout  & ((!\Add0~1 ) # (!\Mux30~1_combout ))))

	.dataa(Mux94),
	.datab(Mux30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~1 ),
	.combout(\Add0~2_combout ),
	.cout(\Add0~3 ));
// synopsys translate_off
defparam \Add0~2 .lut_mask = 16'h9617;
defparam \Add0~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N0
cycloneive_lcell_comb \aluif.portOut[1]~10 (
// Equation(s):
// \aluif.portOut[1]~10_combout  = (\prif.ALUOP_ex [2] & ((\aluif.portOut[1]~9_combout  & (\aluif.portOut[1]~8_combout )) # (!\aluif.portOut[1]~9_combout  & ((\Add0~2_combout ))))) # (!\prif.ALUOP_ex [2] & (\aluif.portOut[1]~9_combout ))

	.dataa(prifALUOP_ex_2),
	.datab(\aluif.portOut[1]~9_combout ),
	.datac(\aluif.portOut[1]~8_combout ),
	.datad(\Add0~2_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[1]~10_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[1]~10 .lut_mask = 16'hE6C4;
defparam \aluif.portOut[1]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N4
cycloneive_lcell_comb \ShiftRight0~6 (
// Equation(s):
// \ShiftRight0~6_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux29~1_combout )) # (!\Mux95~1_combout  & ((\Mux30~1_combout )))))

	.dataa(Mux29),
	.datab(Mux94),
	.datac(Mux30),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~6_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~6 .lut_mask = 16'h2230;
defparam \ShiftRight0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N18
cycloneive_lcell_comb \ShiftRight0~8 (
// Equation(s):
// \ShiftRight0~8_combout  = (!\Mux93~2_combout  & ((\ShiftRight0~6_combout ) # ((\ShiftRight0~7_combout  & \Mux94~1_combout ))))

	.dataa(\ShiftRight0~7_combout ),
	.datab(Mux931),
	.datac(Mux94),
	.datad(\ShiftRight0~6_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~8_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~8 .lut_mask = 16'h3320;
defparam \ShiftRight0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N0
cycloneive_lcell_comb \ShiftRight0~12 (
// Equation(s):
// \ShiftRight0~12_combout  = (!\Mux92~2_combout  & ((\ShiftRight0~8_combout ) # ((\ShiftRight0~11_combout  & \Mux93~2_combout ))))

	.dataa(\ShiftRight0~11_combout ),
	.datab(Mux92),
	.datac(Mux931),
	.datad(\ShiftRight0~8_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~12_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~12 .lut_mask = 16'h3320;
defparam \ShiftRight0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N4
cycloneive_lcell_comb \ShiftRight0~20 (
// Equation(s):
// \ShiftRight0~20_combout  = (!\Mux91~2_combout  & ((\ShiftRight0~12_combout ) # ((\ShiftRight0~19_combout  & \Mux92~2_combout ))))

	.dataa(\ShiftRight0~19_combout ),
	.datab(Mux92),
	.datac(Mux91),
	.datad(\ShiftRight0~12_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~20 .lut_mask = 16'h0F08;
defparam \ShiftRight0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N20
cycloneive_lcell_comb \ShiftRight0~26 (
// Equation(s):
// \ShiftRight0~26_combout  = (\Mux94~1_combout  & (\Mux0~1_combout  & (!\Mux95~1_combout ))) # (!\Mux94~1_combout  & (((\Mux95~1_combout  & \Mux1~1_combout ))))

	.dataa(Mux0),
	.datab(Mux94),
	.datac(Mux95),
	.datad(Mux1),
	.cin(gnd),
	.combout(\ShiftRight0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~26 .lut_mask = 16'h3808;
defparam \ShiftRight0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N18
cycloneive_lcell_comb \ShiftLeft0~16 (
// Equation(s):
// \ShiftLeft0~16_combout  = (!\Mux95~1_combout  & !\Mux94~1_combout )

	.dataa(gnd),
	.datab(Mux95),
	.datac(Mux94),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftLeft0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~16 .lut_mask = 16'h0303;
defparam \ShiftLeft0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N28
cycloneive_lcell_comb \ShiftRight0~27 (
// Equation(s):
// \ShiftRight0~27_combout  = (\Mux93~2_combout  & ((\ShiftRight0~26_combout ) # ((\Mux2~1_combout  & \ShiftLeft0~16_combout ))))

	.dataa(Mux2),
	.datab(\ShiftRight0~26_combout ),
	.datac(Mux931),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~27_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~27 .lut_mask = 16'hE0C0;
defparam \ShiftRight0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N16
cycloneive_lcell_comb \ShiftRight0~22 (
// Equation(s):
// \ShiftRight0~22_combout  = (\ShiftRight0~21_combout  & ((\Mux94~1_combout ) # ((\Mux13~1_combout )))) # (!\ShiftRight0~21_combout  & (!\Mux94~1_combout  & (\Mux14~1_combout )))

	.dataa(\ShiftRight0~21_combout ),
	.datab(Mux94),
	.datac(Mux14),
	.datad(Mux13),
	.cin(gnd),
	.combout(\ShiftRight0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~22 .lut_mask = 16'hBA98;
defparam \ShiftRight0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N24
cycloneive_lcell_comb \ShiftRight0~23 (
// Equation(s):
// \ShiftRight0~23_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux9~1_combout )) # (!\Mux95~1_combout  & ((\Mux10~1_combout )))))

	.dataa(Mux9),
	.datab(Mux95),
	.datac(Mux10),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftRight0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~23 .lut_mask = 16'h00B8;
defparam \ShiftRight0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N22
cycloneive_lcell_comb \ShiftRight0~25 (
// Equation(s):
// \ShiftRight0~25_combout  = (\Mux93~2_combout  & ((\ShiftRight0~24_combout ) # ((\ShiftRight0~23_combout )))) # (!\Mux93~2_combout  & (((\ShiftRight0~22_combout ))))

	.dataa(\ShiftRight0~24_combout ),
	.datab(\ShiftRight0~22_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~23_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~25 .lut_mask = 16'hFCAC;
defparam \ShiftRight0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N26
cycloneive_lcell_comb \ShiftRight0~28 (
// Equation(s):
// \ShiftRight0~28_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux5~1_combout )) # (!\Mux95~1_combout  & ((\Mux6~1_combout )))))

	.dataa(Mux94),
	.datab(Mux5),
	.datac(Mux95),
	.datad(Mux6),
	.cin(gnd),
	.combout(\ShiftRight0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~28 .lut_mask = 16'h4540;
defparam \ShiftRight0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N2
cycloneive_lcell_comb \ShiftRight0~29 (
// Equation(s):
// \ShiftRight0~29_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux3~1_combout ))) # (!\Mux95~1_combout  & (\Mux4~1_combout ))))

	.dataa(Mux94),
	.datab(Mux4),
	.datac(Mux95),
	.datad(Mux3),
	.cin(gnd),
	.combout(\ShiftRight0~29_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~29 .lut_mask = 16'hA808;
defparam \ShiftRight0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N16
cycloneive_lcell_comb \ShiftRight0~30 (
// Equation(s):
// \ShiftRight0~30_combout  = (!\Mux93~2_combout  & ((\ShiftRight0~28_combout ) # (\ShiftRight0~29_combout )))

	.dataa(Mux931),
	.datab(gnd),
	.datac(\ShiftRight0~28_combout ),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~30 .lut_mask = 16'h5550;
defparam \ShiftRight0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N6
cycloneive_lcell_comb \ShiftRight0~31 (
// Equation(s):
// \ShiftRight0~31_combout  = (\Mux92~2_combout  & ((\ShiftRight0~27_combout ) # ((\ShiftRight0~30_combout )))) # (!\Mux92~2_combout  & (((\ShiftRight0~25_combout ))))

	.dataa(Mux92),
	.datab(\ShiftRight0~27_combout ),
	.datac(\ShiftRight0~25_combout ),
	.datad(\ShiftRight0~30_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~31 .lut_mask = 16'hFAD8;
defparam \ShiftRight0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N6
cycloneive_lcell_comb \ShiftRight0~32 (
// Equation(s):
// \ShiftRight0~32_combout  = (\ShiftRight0~20_combout ) # ((\Mux91~2_combout  & \ShiftRight0~31_combout ))

	.dataa(Mux91),
	.datab(gnd),
	.datac(\ShiftRight0~20_combout ),
	.datad(\ShiftRight0~31_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~32 .lut_mask = 16'hFAF0;
defparam \ShiftRight0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N28
cycloneive_lcell_comb \aluif.portOut[1]~13 (
// Equation(s):
// \aluif.portOut[1]~13_combout  = (\prif.ALUOP_ex [2] & \prif.ALUOP_ex [1])

	.dataa(prifALUOP_ex_2),
	.datab(gnd),
	.datac(prifALUOP_ex_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\aluif.portOut[1]~13_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[1]~13 .lut_mask = 16'hA0A0;
defparam \aluif.portOut[1]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N0
cycloneive_lcell_comb \Add1~0 (
// Equation(s):
// \Add1~0_combout  = (\Mux31~1_combout  & ((GND) # (!\Mux95~1_combout ))) # (!\Mux31~1_combout  & (\Mux95~1_combout  $ (GND)))
// \Add1~1  = CARRY((\Mux31~1_combout ) # (!\Mux95~1_combout ))

	.dataa(Mux31),
	.datab(Mux95),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h66BB;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N2
cycloneive_lcell_comb \Add1~2 (
// Equation(s):
// \Add1~2_combout  = (\Mux94~1_combout  & ((\Mux30~1_combout  & (!\Add1~1 )) # (!\Mux30~1_combout  & ((\Add1~1 ) # (GND))))) # (!\Mux94~1_combout  & ((\Mux30~1_combout  & (\Add1~1  & VCC)) # (!\Mux30~1_combout  & (!\Add1~1 ))))
// \Add1~3  = CARRY((\Mux94~1_combout  & ((!\Add1~1 ) # (!\Mux30~1_combout ))) # (!\Mux94~1_combout  & (!\Mux30~1_combout  & !\Add1~1 )))

	.dataa(Mux94),
	.datab(Mux30),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h692B;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N10
cycloneive_lcell_comb \aluif.portOut[1]~11 (
// Equation(s):
// \aluif.portOut[1]~11_combout  = (!\Mux94~1_combout  & !\Mux30~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux94),
	.datad(Mux30),
	.cin(gnd),
	.combout(\aluif.portOut[1]~11_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[1]~11 .lut_mask = 16'h000F;
defparam \aluif.portOut[1]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N4
cycloneive_lcell_comb \aluif.portOut[1]~12 (
// Equation(s):
// \aluif.portOut[1]~12_combout  = (\prif.ALUOP_ex [2] & (!\prif.ALUOP_ex [1] & (\Add1~2_combout ))) # (!\prif.ALUOP_ex [2] & (\prif.ALUOP_ex [1] $ (((\aluif.portOut[1]~11_combout )))))

	.dataa(prifALUOP_ex_2),
	.datab(prifALUOP_ex_1),
	.datac(\Add1~2_combout ),
	.datad(\aluif.portOut[1]~11_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[1]~12_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[1]~12 .lut_mask = 16'h3164;
defparam \aluif.portOut[1]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N28
cycloneive_lcell_comb \aluif.portOut[1]~14 (
// Equation(s):
// \aluif.portOut[1]~14_combout  = (\aluif.portOut[1]~12_combout ) # ((\ShiftRight0~32_combout  & (\aluif.portOut[1]~13_combout  & !\ShiftLeft0~15_combout )))

	.dataa(\ShiftRight0~32_combout ),
	.datab(\aluif.portOut[1]~13_combout ),
	.datac(\aluif.portOut[1]~12_combout ),
	.datad(\ShiftLeft0~15_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[1]~14_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[1]~14 .lut_mask = 16'hF0F8;
defparam \aluif.portOut[1]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N24
cycloneive_lcell_comb \aluif.portOut[0]~16 (
// Equation(s):
// \aluif.portOut[0]~16_combout  = (\prif.ALUOP_ex [2] & (((!\Add1~0_combout )))) # (!\prif.ALUOP_ex [2] & ((\Mux31~1_combout ) # ((\Mux95~1_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(Mux31),
	.datac(Mux95),
	.datad(\Add1~0_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[0]~16_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[0]~16 .lut_mask = 16'h54FE;
defparam \aluif.portOut[0]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N8
cycloneive_lcell_comb \aluif.portOut[0]~17 (
// Equation(s):
// \aluif.portOut[0]~17_combout  = (\prif.ALUOP_ex [0] & (\Add0~0_combout )) # (!\prif.ALUOP_ex [0] & ((!\aluif.portOut[0]~16_combout )))

	.dataa(\Add0~0_combout ),
	.datab(prifALUOP_ex_0),
	.datac(gnd),
	.datad(\aluif.portOut[0]~16_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[0]~17_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[0]~17 .lut_mask = 16'h88BB;
defparam \aluif.portOut[0]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N4
cycloneive_lcell_comb \ShiftRight0~53 (
// Equation(s):
// \ShiftRight0~53_combout  = (\Mux95~1_combout  & ((\Mux16~1_combout ))) # (!\Mux95~1_combout  & (\Mux17~1_combout ))

	.dataa(gnd),
	.datab(Mux17),
	.datac(Mux95),
	.datad(Mux16),
	.cin(gnd),
	.combout(\ShiftRight0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~53 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N6
cycloneive_lcell_comb \ShiftRight0~54 (
// Equation(s):
// \ShiftRight0~54_combout  = (\Mux95~1_combout  & (((\Mux18~1_combout )))) # (!\Mux95~1_combout  & ((\Mux19~1_combout ) # ((\Mux19~0_combout ))))

	.dataa(Mux191),
	.datab(Mux19),
	.datac(Mux18),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~54 .lut_mask = 16'hF0EE;
defparam \ShiftRight0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N22
cycloneive_lcell_comb \ShiftRight0~55 (
// Equation(s):
// \ShiftRight0~55_combout  = (\Mux94~1_combout  & (\ShiftRight0~53_combout )) # (!\Mux94~1_combout  & ((\ShiftRight0~54_combout )))

	.dataa(Mux94),
	.datab(gnd),
	.datac(\ShiftRight0~53_combout ),
	.datad(\ShiftRight0~54_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~55 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N18
cycloneive_lcell_comb \ShiftRight0~57 (
// Equation(s):
// \ShiftRight0~57_combout  = (\Mux95~1_combout  & (\Mux22~1_combout )) # (!\Mux95~1_combout  & ((\Mux23~1_combout )))

	.dataa(gnd),
	.datab(Mux22),
	.datac(Mux95),
	.datad(Mux23),
	.cin(gnd),
	.combout(\ShiftRight0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~57 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N20
cycloneive_lcell_comb \ShiftRight0~56 (
// Equation(s):
// \ShiftRight0~56_combout  = (\Mux95~1_combout  & (\Mux20~1_combout )) # (!\Mux95~1_combout  & ((\Mux21~1_combout )))

	.dataa(gnd),
	.datab(Mux95),
	.datac(Mux20),
	.datad(Mux21),
	.cin(gnd),
	.combout(\ShiftRight0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~56 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N28
cycloneive_lcell_comb \ShiftRight0~58 (
// Equation(s):
// \ShiftRight0~58_combout  = (\Mux94~1_combout  & ((\ShiftRight0~56_combout ))) # (!\Mux94~1_combout  & (\ShiftRight0~57_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~57_combout ),
	.datac(Mux94),
	.datad(\ShiftRight0~56_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~58 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N10
cycloneive_lcell_comb \ShiftRight0~59 (
// Equation(s):
// \ShiftRight0~59_combout  = (\Mux93~2_combout  & (\ShiftRight0~55_combout )) # (!\Mux93~2_combout  & ((\ShiftRight0~58_combout )))

	.dataa(gnd),
	.datab(Mux931),
	.datac(\ShiftRight0~55_combout ),
	.datad(\ShiftRight0~58_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~59 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N8
cycloneive_lcell_comb \ShiftRight0~50 (
// Equation(s):
// \ShiftRight0~50_combout  = (\Mux95~1_combout  & (\Mux26~1_combout )) # (!\Mux95~1_combout  & ((\Mux27~1_combout )))

	.dataa(gnd),
	.datab(Mux95),
	.datac(Mux26),
	.datad(Mux27),
	.cin(gnd),
	.combout(\ShiftRight0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~50 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N30
cycloneive_lcell_comb \ShiftRight0~49 (
// Equation(s):
// \ShiftRight0~49_combout  = (\Mux95~1_combout  & (\Mux24~1_combout )) # (!\Mux95~1_combout  & ((\Mux25~1_combout )))

	.dataa(Mux24),
	.datab(Mux95),
	.datac(gnd),
	.datad(Mux25),
	.cin(gnd),
	.combout(\ShiftRight0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~49 .lut_mask = 16'hBB88;
defparam \ShiftRight0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N22
cycloneive_lcell_comb \ShiftRight0~51 (
// Equation(s):
// \ShiftRight0~51_combout  = (\Mux94~1_combout  & ((\ShiftRight0~49_combout ))) # (!\Mux94~1_combout  & (\ShiftRight0~50_combout ))

	.dataa(Mux94),
	.datab(\ShiftRight0~50_combout ),
	.datac(\ShiftRight0~49_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~51 .lut_mask = 16'hE4E4;
defparam \ShiftRight0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N14
cycloneive_lcell_comb \ShiftRight0~47 (
// Equation(s):
// \ShiftRight0~47_combout  = (\Mux95~1_combout  & ((\Mux28~1_combout ))) # (!\Mux95~1_combout  & (\Mux29~1_combout ))

	.dataa(Mux29),
	.datab(Mux95),
	.datac(gnd),
	.datad(Mux28),
	.cin(gnd),
	.combout(\ShiftRight0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~47 .lut_mask = 16'hEE22;
defparam \ShiftRight0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N0
cycloneive_lcell_comb \ShiftRight0~48 (
// Equation(s):
// \ShiftRight0~48_combout  = (!\Mux93~2_combout  & ((\ShiftRight0~46_combout ) # ((\Mux94~1_combout  & \ShiftRight0~47_combout ))))

	.dataa(\ShiftRight0~46_combout ),
	.datab(Mux931),
	.datac(Mux94),
	.datad(\ShiftRight0~47_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~48 .lut_mask = 16'h3222;
defparam \ShiftRight0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N20
cycloneive_lcell_comb \ShiftRight0~52 (
// Equation(s):
// \ShiftRight0~52_combout  = (!\Mux92~2_combout  & ((\ShiftRight0~48_combout ) # ((\Mux93~2_combout  & \ShiftRight0~51_combout ))))

	.dataa(Mux92),
	.datab(Mux931),
	.datac(\ShiftRight0~51_combout ),
	.datad(\ShiftRight0~48_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~52_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~52 .lut_mask = 16'h5540;
defparam \ShiftRight0~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N8
cycloneive_lcell_comb \ShiftRight0~60 (
// Equation(s):
// \ShiftRight0~60_combout  = (\ShiftRight0~52_combout ) # ((\Mux92~2_combout  & \ShiftRight0~59_combout ))

	.dataa(Mux92),
	.datab(gnd),
	.datac(\ShiftRight0~59_combout ),
	.datad(\ShiftRight0~52_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~60 .lut_mask = 16'hFFA0;
defparam \ShiftRight0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N2
cycloneive_lcell_comb \aluif.portOut[0]~18 (
// Equation(s):
// \aluif.portOut[0]~18_combout  = ((\Mux91~2_combout  & (\ShiftRight0~45_combout )) # (!\Mux91~2_combout  & ((\ShiftRight0~60_combout )))) # (!\prif.ALUOP_ex [2])

	.dataa(\ShiftRight0~45_combout ),
	.datab(\ShiftRight0~60_combout ),
	.datac(prifALUOP_ex_2),
	.datad(Mux91),
	.cin(gnd),
	.combout(\aluif.portOut[0]~18_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[0]~18 .lut_mask = 16'hAFCF;
defparam \aluif.portOut[0]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N22
cycloneive_lcell_comb \portOut~1 (
// Equation(s):
// \portOut~1_combout  = (\Mux95~1_combout ) # (\Mux31~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux95),
	.datad(Mux31),
	.cin(gnd),
	.combout(\portOut~1_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~1 .lut_mask = 16'hFFF0;
defparam \portOut~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N18
cycloneive_lcell_comb \aluif.portOut[0]~20 (
// Equation(s):
// \aluif.portOut[0]~20_combout  = (\prif.ALUOP_ex [2] & (\prif.ALUOP_ex [0] $ ((!\ShiftLeft0~15_combout )))) # (!\prif.ALUOP_ex [2] & (!\prif.ALUOP_ex [0] & ((\portOut~1_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(prifALUOP_ex_0),
	.datac(\ShiftLeft0~15_combout ),
	.datad(\portOut~1_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[0]~20_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[0]~20 .lut_mask = 16'h9382;
defparam \aluif.portOut[0]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N12
cycloneive_lcell_comb \aluif.portOut[0]~21 (
// Equation(s):
// \aluif.portOut[0]~21_combout  = (\prif.ALUOP_ex [0] & (\aluif.portOut[0]~19_combout  & ((!\aluif.portOut[0]~20_combout )))) # (!\prif.ALUOP_ex [0] & (((\aluif.portOut[0]~18_combout  & \aluif.portOut[0]~20_combout ))))

	.dataa(\aluif.portOut[0]~19_combout ),
	.datab(prifALUOP_ex_0),
	.datac(\aluif.portOut[0]~18_combout ),
	.datad(\aluif.portOut[0]~20_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[0]~21_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[0]~21 .lut_mask = 16'h3088;
defparam \aluif.portOut[0]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N30
cycloneive_lcell_comb \aluif.portOut[0]~22 (
// Equation(s):
// \aluif.portOut[0]~22_combout  = (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [1] & ((\aluif.portOut[0]~21_combout ))) # (!\prif.ALUOP_ex [1] & (\aluif.portOut[0]~17_combout ))))

	.dataa(prifALUOP_ex_1),
	.datab(\aluif.portOut[0]~17_combout ),
	.datac(prifALUOP_ex_3),
	.datad(\aluif.portOut[0]~21_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[0]~22_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[0]~22 .lut_mask = 16'hE040;
defparam \aluif.portOut[0]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N0
cycloneive_lcell_comb \LessThan0~1 (
// Equation(s):
// \LessThan0~1_cout  = CARRY((\Mux95~1_combout  & !\Mux31~1_combout ))

	.dataa(Mux95),
	.datab(Mux31),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan0~1_cout ));
// synopsys translate_off
defparam \LessThan0~1 .lut_mask = 16'h0022;
defparam \LessThan0~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N2
cycloneive_lcell_comb \LessThan0~3 (
// Equation(s):
// \LessThan0~3_cout  = CARRY((\Mux94~1_combout  & (\Mux30~1_combout  & !\LessThan0~1_cout )) # (!\Mux94~1_combout  & ((\Mux30~1_combout ) # (!\LessThan0~1_cout ))))

	.dataa(Mux94),
	.datab(Mux30),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~1_cout ),
	.combout(),
	.cout(\LessThan0~3_cout ));
// synopsys translate_off
defparam \LessThan0~3 .lut_mask = 16'h004D;
defparam \LessThan0~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N4
cycloneive_lcell_comb \LessThan0~5 (
// Equation(s):
// \LessThan0~5_cout  = CARRY((\Mux93~2_combout  & ((!\LessThan0~3_cout ) # (!\Mux29~1_combout ))) # (!\Mux93~2_combout  & (!\Mux29~1_combout  & !\LessThan0~3_cout )))

	.dataa(Mux931),
	.datab(Mux29),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~3_cout ),
	.combout(),
	.cout(\LessThan0~5_cout ));
// synopsys translate_off
defparam \LessThan0~5 .lut_mask = 16'h002B;
defparam \LessThan0~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N6
cycloneive_lcell_comb \LessThan0~7 (
// Equation(s):
// \LessThan0~7_cout  = CARRY((\Mux92~2_combout  & (\Mux28~1_combout  & !\LessThan0~5_cout )) # (!\Mux92~2_combout  & ((\Mux28~1_combout ) # (!\LessThan0~5_cout ))))

	.dataa(Mux92),
	.datab(Mux28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~5_cout ),
	.combout(),
	.cout(\LessThan0~7_cout ));
// synopsys translate_off
defparam \LessThan0~7 .lut_mask = 16'h004D;
defparam \LessThan0~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N8
cycloneive_lcell_comb \LessThan0~9 (
// Equation(s):
// \LessThan0~9_cout  = CARRY((\Mux91~2_combout  & ((!\LessThan0~7_cout ) # (!\Mux27~1_combout ))) # (!\Mux91~2_combout  & (!\Mux27~1_combout  & !\LessThan0~7_cout )))

	.dataa(Mux91),
	.datab(Mux27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~7_cout ),
	.combout(),
	.cout(\LessThan0~9_cout ));
// synopsys translate_off
defparam \LessThan0~9 .lut_mask = 16'h002B;
defparam \LessThan0~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N10
cycloneive_lcell_comb \LessThan0~11 (
// Equation(s):
// \LessThan0~11_cout  = CARRY((\Mux90~3_combout  & (\Mux26~1_combout  & !\LessThan0~9_cout )) # (!\Mux90~3_combout  & ((\Mux26~1_combout ) # (!\LessThan0~9_cout ))))

	.dataa(Mux90),
	.datab(Mux26),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~9_cout ),
	.combout(),
	.cout(\LessThan0~11_cout ));
// synopsys translate_off
defparam \LessThan0~11 .lut_mask = 16'h004D;
defparam \LessThan0~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N12
cycloneive_lcell_comb \LessThan0~13 (
// Equation(s):
// \LessThan0~13_cout  = CARRY((\Mux89~4_combout  & ((!\LessThan0~11_cout ) # (!\Mux25~1_combout ))) # (!\Mux89~4_combout  & (!\Mux25~1_combout  & !\LessThan0~11_cout )))

	.dataa(Mux891),
	.datab(Mux25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~11_cout ),
	.combout(),
	.cout(\LessThan0~13_cout ));
// synopsys translate_off
defparam \LessThan0~13 .lut_mask = 16'h002B;
defparam \LessThan0~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N14
cycloneive_lcell_comb \LessThan0~15 (
// Equation(s):
// \LessThan0~15_cout  = CARRY((\Mux88~3_combout  & (\Mux24~1_combout  & !\LessThan0~13_cout )) # (!\Mux88~3_combout  & ((\Mux24~1_combout ) # (!\LessThan0~13_cout ))))

	.dataa(Mux88),
	.datab(Mux24),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~13_cout ),
	.combout(),
	.cout(\LessThan0~15_cout ));
// synopsys translate_off
defparam \LessThan0~15 .lut_mask = 16'h004D;
defparam \LessThan0~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N16
cycloneive_lcell_comb \LessThan0~17 (
// Equation(s):
// \LessThan0~17_cout  = CARRY((\Mux23~1_combout  & (\Mux87~3_combout  & !\LessThan0~15_cout )) # (!\Mux23~1_combout  & ((\Mux87~3_combout ) # (!\LessThan0~15_cout ))))

	.dataa(Mux23),
	.datab(Mux87),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~15_cout ),
	.combout(),
	.cout(\LessThan0~17_cout ));
// synopsys translate_off
defparam \LessThan0~17 .lut_mask = 16'h004D;
defparam \LessThan0~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N18
cycloneive_lcell_comb \LessThan0~19 (
// Equation(s):
// \LessThan0~19_cout  = CARRY((\Mux22~1_combout  & ((!\LessThan0~17_cout ) # (!\Mux86~3_combout ))) # (!\Mux22~1_combout  & (!\Mux86~3_combout  & !\LessThan0~17_cout )))

	.dataa(Mux22),
	.datab(Mux86),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~17_cout ),
	.combout(),
	.cout(\LessThan0~19_cout ));
// synopsys translate_off
defparam \LessThan0~19 .lut_mask = 16'h002B;
defparam \LessThan0~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N20
cycloneive_lcell_comb \LessThan0~21 (
// Equation(s):
// \LessThan0~21_cout  = CARRY((\Mux85~3_combout  & ((!\LessThan0~19_cout ) # (!\Mux21~1_combout ))) # (!\Mux85~3_combout  & (!\Mux21~1_combout  & !\LessThan0~19_cout )))

	.dataa(Mux85),
	.datab(Mux21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~19_cout ),
	.combout(),
	.cout(\LessThan0~21_cout ));
// synopsys translate_off
defparam \LessThan0~21 .lut_mask = 16'h002B;
defparam \LessThan0~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N22
cycloneive_lcell_comb \LessThan0~23 (
// Equation(s):
// \LessThan0~23_cout  = CARRY((\Mux84~3_combout  & (\Mux20~1_combout  & !\LessThan0~21_cout )) # (!\Mux84~3_combout  & ((\Mux20~1_combout ) # (!\LessThan0~21_cout ))))

	.dataa(Mux84),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~21_cout ),
	.combout(),
	.cout(\LessThan0~23_cout ));
// synopsys translate_off
defparam \LessThan0~23 .lut_mask = 16'h004D;
defparam \LessThan0~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N24
cycloneive_lcell_comb \LessThan0~25 (
// Equation(s):
// \LessThan0~25_cout  = CARRY((\Mux19~3_combout  & (\Mux83~3_combout  & !\LessThan0~23_cout )) # (!\Mux19~3_combout  & ((\Mux83~3_combout ) # (!\LessThan0~23_cout ))))

	.dataa(Mux192),
	.datab(Mux83),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~23_cout ),
	.combout(),
	.cout(\LessThan0~25_cout ));
// synopsys translate_off
defparam \LessThan0~25 .lut_mask = 16'h004D;
defparam \LessThan0~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N26
cycloneive_lcell_comb \LessThan0~27 (
// Equation(s):
// \LessThan0~27_cout  = CARRY((\Mux82~3_combout  & (\Mux18~1_combout  & !\LessThan0~25_cout )) # (!\Mux82~3_combout  & ((\Mux18~1_combout ) # (!\LessThan0~25_cout ))))

	.dataa(Mux82),
	.datab(Mux18),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~25_cout ),
	.combout(),
	.cout(\LessThan0~27_cout ));
// synopsys translate_off
defparam \LessThan0~27 .lut_mask = 16'h004D;
defparam \LessThan0~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N28
cycloneive_lcell_comb \LessThan0~29 (
// Equation(s):
// \LessThan0~29_cout  = CARRY((\Mux17~1_combout  & (\Mux81~3_combout  & !\LessThan0~27_cout )) # (!\Mux17~1_combout  & ((\Mux81~3_combout ) # (!\LessThan0~27_cout ))))

	.dataa(Mux17),
	.datab(Mux81),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~27_cout ),
	.combout(),
	.cout(\LessThan0~29_cout ));
// synopsys translate_off
defparam \LessThan0~29 .lut_mask = 16'h004D;
defparam \LessThan0~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y26_N30
cycloneive_lcell_comb \LessThan0~31 (
// Equation(s):
// \LessThan0~31_cout  = CARRY((\Mux80~4_combout  & (\Mux16~1_combout  & !\LessThan0~29_cout )) # (!\Mux80~4_combout  & ((\Mux16~1_combout ) # (!\LessThan0~29_cout ))))

	.dataa(Mux80),
	.datab(Mux16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~29_cout ),
	.combout(),
	.cout(\LessThan0~31_cout ));
// synopsys translate_off
defparam \LessThan0~31 .lut_mask = 16'h004D;
defparam \LessThan0~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N0
cycloneive_lcell_comb \LessThan0~33 (
// Equation(s):
// \LessThan0~33_cout  = CARRY((\Mux79~0_combout  & ((!\LessThan0~31_cout ) # (!\Mux15~1_combout ))) # (!\Mux79~0_combout  & (!\Mux15~1_combout  & !\LessThan0~31_cout )))

	.dataa(Mux79),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~31_cout ),
	.combout(),
	.cout(\LessThan0~33_cout ));
// synopsys translate_off
defparam \LessThan0~33 .lut_mask = 16'h002B;
defparam \LessThan0~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N2
cycloneive_lcell_comb \LessThan0~35 (
// Equation(s):
// \LessThan0~35_cout  = CARRY((\Mux14~1_combout  & ((!\LessThan0~33_cout ) # (!\Mux78~0_combout ))) # (!\Mux14~1_combout  & (!\Mux78~0_combout  & !\LessThan0~33_cout )))

	.dataa(Mux14),
	.datab(Mux78),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~33_cout ),
	.combout(),
	.cout(\LessThan0~35_cout ));
// synopsys translate_off
defparam \LessThan0~35 .lut_mask = 16'h002B;
defparam \LessThan0~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N4
cycloneive_lcell_comb \LessThan0~37 (
// Equation(s):
// \LessThan0~37_cout  = CARRY((\Mux77~0_combout  & ((!\LessThan0~35_cout ) # (!\Mux13~1_combout ))) # (!\Mux77~0_combout  & (!\Mux13~1_combout  & !\LessThan0~35_cout )))

	.dataa(Mux77),
	.datab(Mux13),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~35_cout ),
	.combout(),
	.cout(\LessThan0~37_cout ));
// synopsys translate_off
defparam \LessThan0~37 .lut_mask = 16'h002B;
defparam \LessThan0~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N6
cycloneive_lcell_comb \LessThan0~39 (
// Equation(s):
// \LessThan0~39_cout  = CARRY((\Mux12~1_combout  & ((!\LessThan0~37_cout ) # (!\Mux76~0_combout ))) # (!\Mux12~1_combout  & (!\Mux76~0_combout  & !\LessThan0~37_cout )))

	.dataa(Mux12),
	.datab(Mux76),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~37_cout ),
	.combout(),
	.cout(\LessThan0~39_cout ));
// synopsys translate_off
defparam \LessThan0~39 .lut_mask = 16'h002B;
defparam \LessThan0~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N8
cycloneive_lcell_comb \LessThan0~41 (
// Equation(s):
// \LessThan0~41_cout  = CARRY((\Mux11~1_combout  & (\Mux75~0_combout  & !\LessThan0~39_cout )) # (!\Mux11~1_combout  & ((\Mux75~0_combout ) # (!\LessThan0~39_cout ))))

	.dataa(Mux11),
	.datab(Mux75),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~39_cout ),
	.combout(),
	.cout(\LessThan0~41_cout ));
// synopsys translate_off
defparam \LessThan0~41 .lut_mask = 16'h004D;
defparam \LessThan0~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N10
cycloneive_lcell_comb \LessThan0~43 (
// Equation(s):
// \LessThan0~43_cout  = CARRY((\Mux74~0_combout  & (\Mux10~1_combout  & !\LessThan0~41_cout )) # (!\Mux74~0_combout  & ((\Mux10~1_combout ) # (!\LessThan0~41_cout ))))

	.dataa(Mux74),
	.datab(Mux10),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~41_cout ),
	.combout(),
	.cout(\LessThan0~43_cout ));
// synopsys translate_off
defparam \LessThan0~43 .lut_mask = 16'h004D;
defparam \LessThan0~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N12
cycloneive_lcell_comb \LessThan0~45 (
// Equation(s):
// \LessThan0~45_cout  = CARRY((\Mux9~1_combout  & (\Mux73~0_combout  & !\LessThan0~43_cout )) # (!\Mux9~1_combout  & ((\Mux73~0_combout ) # (!\LessThan0~43_cout ))))

	.dataa(Mux9),
	.datab(Mux73),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~43_cout ),
	.combout(),
	.cout(\LessThan0~45_cout ));
// synopsys translate_off
defparam \LessThan0~45 .lut_mask = 16'h004D;
defparam \LessThan0~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N14
cycloneive_lcell_comb \LessThan0~47 (
// Equation(s):
// \LessThan0~47_cout  = CARRY((\Mux8~1_combout  & ((!\LessThan0~45_cout ) # (!\Mux72~0_combout ))) # (!\Mux8~1_combout  & (!\Mux72~0_combout  & !\LessThan0~45_cout )))

	.dataa(Mux8),
	.datab(Mux72),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~45_cout ),
	.combout(),
	.cout(\LessThan0~47_cout ));
// synopsys translate_off
defparam \LessThan0~47 .lut_mask = 16'h002B;
defparam \LessThan0~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N16
cycloneive_lcell_comb \LessThan0~49 (
// Equation(s):
// \LessThan0~49_cout  = CARRY((\Mux71~0_combout  & ((!\LessThan0~47_cout ) # (!\Mux7~1_combout ))) # (!\Mux71~0_combout  & (!\Mux7~1_combout  & !\LessThan0~47_cout )))

	.dataa(Mux71),
	.datab(Mux7),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~47_cout ),
	.combout(),
	.cout(\LessThan0~49_cout ));
// synopsys translate_off
defparam \LessThan0~49 .lut_mask = 16'h002B;
defparam \LessThan0~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N18
cycloneive_lcell_comb \LessThan0~51 (
// Equation(s):
// \LessThan0~51_cout  = CARRY((\Mux6~1_combout  & ((!\LessThan0~49_cout ) # (!\Mux70~0_combout ))) # (!\Mux6~1_combout  & (!\Mux70~0_combout  & !\LessThan0~49_cout )))

	.dataa(Mux6),
	.datab(Mux70),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~49_cout ),
	.combout(),
	.cout(\LessThan0~51_cout ));
// synopsys translate_off
defparam \LessThan0~51 .lut_mask = 16'h002B;
defparam \LessThan0~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N20
cycloneive_lcell_comb \LessThan0~53 (
// Equation(s):
// \LessThan0~53_cout  = CARRY((\Mux69~0_combout  & ((!\LessThan0~51_cout ) # (!\Mux5~1_combout ))) # (!\Mux69~0_combout  & (!\Mux5~1_combout  & !\LessThan0~51_cout )))

	.dataa(Mux69),
	.datab(Mux5),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~51_cout ),
	.combout(),
	.cout(\LessThan0~53_cout ));
// synopsys translate_off
defparam \LessThan0~53 .lut_mask = 16'h002B;
defparam \LessThan0~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N22
cycloneive_lcell_comb \LessThan0~55 (
// Equation(s):
// \LessThan0~55_cout  = CARRY((\Mux68~0_combout  & (\Mux4~1_combout  & !\LessThan0~53_cout )) # (!\Mux68~0_combout  & ((\Mux4~1_combout ) # (!\LessThan0~53_cout ))))

	.dataa(Mux68),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~53_cout ),
	.combout(),
	.cout(\LessThan0~55_cout ));
// synopsys translate_off
defparam \LessThan0~55 .lut_mask = 16'h004D;
defparam \LessThan0~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N24
cycloneive_lcell_comb \LessThan0~57 (
// Equation(s):
// \LessThan0~57_cout  = CARRY((\Mux67~0_combout  & ((!\LessThan0~55_cout ) # (!\Mux3~1_combout ))) # (!\Mux67~0_combout  & (!\Mux3~1_combout  & !\LessThan0~55_cout )))

	.dataa(Mux67),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~55_cout ),
	.combout(),
	.cout(\LessThan0~57_cout ));
// synopsys translate_off
defparam \LessThan0~57 .lut_mask = 16'h002B;
defparam \LessThan0~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N26
cycloneive_lcell_comb \LessThan0~59 (
// Equation(s):
// \LessThan0~59_cout  = CARRY((\Mux66~0_combout  & (\Mux2~1_combout  & !\LessThan0~57_cout )) # (!\Mux66~0_combout  & ((\Mux2~1_combout ) # (!\LessThan0~57_cout ))))

	.dataa(Mux66),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~57_cout ),
	.combout(),
	.cout(\LessThan0~59_cout ));
// synopsys translate_off
defparam \LessThan0~59 .lut_mask = 16'h004D;
defparam \LessThan0~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N28
cycloneive_lcell_comb \LessThan0~61 (
// Equation(s):
// \LessThan0~61_cout  = CARRY((\Mux65~0_combout  & ((!\LessThan0~59_cout ) # (!\Mux1~1_combout ))) # (!\Mux65~0_combout  & (!\Mux1~1_combout  & !\LessThan0~59_cout )))

	.dataa(Mux65),
	.datab(Mux1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan0~59_cout ),
	.combout(),
	.cout(\LessThan0~61_cout ));
// synopsys translate_off
defparam \LessThan0~61 .lut_mask = 16'h002B;
defparam \LessThan0~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y25_N30
cycloneive_lcell_comb \LessThan0~62 (
// Equation(s):
// \LessThan0~62_combout  = (\Mux0~1_combout  & ((\LessThan0~61_cout ) # (!\Mux64~0_combout ))) # (!\Mux0~1_combout  & (\LessThan0~61_cout  & !\Mux64~0_combout ))

	.dataa(Mux0),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux64),
	.cin(\LessThan0~61_cout ),
	.combout(\LessThan0~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan0~62 .lut_mask = 16'hA0FA;
defparam \LessThan0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N0
cycloneive_lcell_comb \LessThan1~1 (
// Equation(s):
// \LessThan1~1_cout  = CARRY((!\Mux31~1_combout  & \Mux95~1_combout ))

	.dataa(Mux31),
	.datab(Mux95),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(),
	.cout(\LessThan1~1_cout ));
// synopsys translate_off
defparam \LessThan1~1 .lut_mask = 16'h0044;
defparam \LessThan1~1 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N2
cycloneive_lcell_comb \LessThan1~3 (
// Equation(s):
// \LessThan1~3_cout  = CARRY((\Mux30~1_combout  & ((!\LessThan1~1_cout ) # (!\Mux94~1_combout ))) # (!\Mux30~1_combout  & (!\Mux94~1_combout  & !\LessThan1~1_cout )))

	.dataa(Mux30),
	.datab(Mux94),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~1_cout ),
	.combout(),
	.cout(\LessThan1~3_cout ));
// synopsys translate_off
defparam \LessThan1~3 .lut_mask = 16'h002B;
defparam \LessThan1~3 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N4
cycloneive_lcell_comb \LessThan1~5 (
// Equation(s):
// \LessThan1~5_cout  = CARRY((\Mux29~1_combout  & (\Mux93~2_combout  & !\LessThan1~3_cout )) # (!\Mux29~1_combout  & ((\Mux93~2_combout ) # (!\LessThan1~3_cout ))))

	.dataa(Mux29),
	.datab(Mux931),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~3_cout ),
	.combout(),
	.cout(\LessThan1~5_cout ));
// synopsys translate_off
defparam \LessThan1~5 .lut_mask = 16'h004D;
defparam \LessThan1~5 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N6
cycloneive_lcell_comb \LessThan1~7 (
// Equation(s):
// \LessThan1~7_cout  = CARRY((\Mux92~2_combout  & (\Mux28~1_combout  & !\LessThan1~5_cout )) # (!\Mux92~2_combout  & ((\Mux28~1_combout ) # (!\LessThan1~5_cout ))))

	.dataa(Mux92),
	.datab(Mux28),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~5_cout ),
	.combout(),
	.cout(\LessThan1~7_cout ));
// synopsys translate_off
defparam \LessThan1~7 .lut_mask = 16'h004D;
defparam \LessThan1~7 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N8
cycloneive_lcell_comb \LessThan1~9 (
// Equation(s):
// \LessThan1~9_cout  = CARRY((\Mux91~2_combout  & ((!\LessThan1~7_cout ) # (!\Mux27~1_combout ))) # (!\Mux91~2_combout  & (!\Mux27~1_combout  & !\LessThan1~7_cout )))

	.dataa(Mux91),
	.datab(Mux27),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~7_cout ),
	.combout(),
	.cout(\LessThan1~9_cout ));
// synopsys translate_off
defparam \LessThan1~9 .lut_mask = 16'h002B;
defparam \LessThan1~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N10
cycloneive_lcell_comb \LessThan1~11 (
// Equation(s):
// \LessThan1~11_cout  = CARRY((\Mux26~1_combout  & ((!\LessThan1~9_cout ) # (!\Mux90~3_combout ))) # (!\Mux26~1_combout  & (!\Mux90~3_combout  & !\LessThan1~9_cout )))

	.dataa(Mux26),
	.datab(Mux90),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~9_cout ),
	.combout(),
	.cout(\LessThan1~11_cout ));
// synopsys translate_off
defparam \LessThan1~11 .lut_mask = 16'h002B;
defparam \LessThan1~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N12
cycloneive_lcell_comb \LessThan1~13 (
// Equation(s):
// \LessThan1~13_cout  = CARRY((\Mux89~4_combout  & ((!\LessThan1~11_cout ) # (!\Mux25~1_combout ))) # (!\Mux89~4_combout  & (!\Mux25~1_combout  & !\LessThan1~11_cout )))

	.dataa(Mux891),
	.datab(Mux25),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~11_cout ),
	.combout(),
	.cout(\LessThan1~13_cout ));
// synopsys translate_off
defparam \LessThan1~13 .lut_mask = 16'h002B;
defparam \LessThan1~13 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N14
cycloneive_lcell_comb \LessThan1~15 (
// Equation(s):
// \LessThan1~15_cout  = CARRY((\Mux24~1_combout  & ((!\LessThan1~13_cout ) # (!\Mux88~3_combout ))) # (!\Mux24~1_combout  & (!\Mux88~3_combout  & !\LessThan1~13_cout )))

	.dataa(Mux24),
	.datab(Mux88),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~13_cout ),
	.combout(),
	.cout(\LessThan1~15_cout ));
// synopsys translate_off
defparam \LessThan1~15 .lut_mask = 16'h002B;
defparam \LessThan1~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N16
cycloneive_lcell_comb \LessThan1~17 (
// Equation(s):
// \LessThan1~17_cout  = CARRY((\Mux23~1_combout  & (\Mux87~3_combout  & !\LessThan1~15_cout )) # (!\Mux23~1_combout  & ((\Mux87~3_combout ) # (!\LessThan1~15_cout ))))

	.dataa(Mux23),
	.datab(Mux87),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~15_cout ),
	.combout(),
	.cout(\LessThan1~17_cout ));
// synopsys translate_off
defparam \LessThan1~17 .lut_mask = 16'h004D;
defparam \LessThan1~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N18
cycloneive_lcell_comb \LessThan1~19 (
// Equation(s):
// \LessThan1~19_cout  = CARRY((\Mux22~1_combout  & ((!\LessThan1~17_cout ) # (!\Mux86~3_combout ))) # (!\Mux22~1_combout  & (!\Mux86~3_combout  & !\LessThan1~17_cout )))

	.dataa(Mux22),
	.datab(Mux86),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~17_cout ),
	.combout(),
	.cout(\LessThan1~19_cout ));
// synopsys translate_off
defparam \LessThan1~19 .lut_mask = 16'h002B;
defparam \LessThan1~19 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N20
cycloneive_lcell_comb \LessThan1~21 (
// Equation(s):
// \LessThan1~21_cout  = CARRY((\Mux85~3_combout  & ((!\LessThan1~19_cout ) # (!\Mux21~1_combout ))) # (!\Mux85~3_combout  & (!\Mux21~1_combout  & !\LessThan1~19_cout )))

	.dataa(Mux85),
	.datab(Mux21),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~19_cout ),
	.combout(),
	.cout(\LessThan1~21_cout ));
// synopsys translate_off
defparam \LessThan1~21 .lut_mask = 16'h002B;
defparam \LessThan1~21 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N22
cycloneive_lcell_comb \LessThan1~23 (
// Equation(s):
// \LessThan1~23_cout  = CARRY((\Mux84~3_combout  & (\Mux20~1_combout  & !\LessThan1~21_cout )) # (!\Mux84~3_combout  & ((\Mux20~1_combout ) # (!\LessThan1~21_cout ))))

	.dataa(Mux84),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~21_cout ),
	.combout(),
	.cout(\LessThan1~23_cout ));
// synopsys translate_off
defparam \LessThan1~23 .lut_mask = 16'h004D;
defparam \LessThan1~23 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N24
cycloneive_lcell_comb \LessThan1~25 (
// Equation(s):
// \LessThan1~25_cout  = CARRY((\Mux83~3_combout  & ((!\LessThan1~23_cout ) # (!\Mux19~3_combout ))) # (!\Mux83~3_combout  & (!\Mux19~3_combout  & !\LessThan1~23_cout )))

	.dataa(Mux83),
	.datab(Mux192),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~23_cout ),
	.combout(),
	.cout(\LessThan1~25_cout ));
// synopsys translate_off
defparam \LessThan1~25 .lut_mask = 16'h002B;
defparam \LessThan1~25 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N26
cycloneive_lcell_comb \LessThan1~27 (
// Equation(s):
// \LessThan1~27_cout  = CARRY((\Mux18~1_combout  & ((!\LessThan1~25_cout ) # (!\Mux82~3_combout ))) # (!\Mux18~1_combout  & (!\Mux82~3_combout  & !\LessThan1~25_cout )))

	.dataa(Mux18),
	.datab(Mux82),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~25_cout ),
	.combout(),
	.cout(\LessThan1~27_cout ));
// synopsys translate_off
defparam \LessThan1~27 .lut_mask = 16'h002B;
defparam \LessThan1~27 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N28
cycloneive_lcell_comb \LessThan1~29 (
// Equation(s):
// \LessThan1~29_cout  = CARRY((\Mux81~3_combout  & ((!\LessThan1~27_cout ) # (!\Mux17~1_combout ))) # (!\Mux81~3_combout  & (!\Mux17~1_combout  & !\LessThan1~27_cout )))

	.dataa(Mux81),
	.datab(Mux17),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~27_cout ),
	.combout(),
	.cout(\LessThan1~29_cout ));
// synopsys translate_off
defparam \LessThan1~29 .lut_mask = 16'h002B;
defparam \LessThan1~29 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y24_N30
cycloneive_lcell_comb \LessThan1~31 (
// Equation(s):
// \LessThan1~31_cout  = CARRY((\Mux80~4_combout  & (\Mux16~1_combout  & !\LessThan1~29_cout )) # (!\Mux80~4_combout  & ((\Mux16~1_combout ) # (!\LessThan1~29_cout ))))

	.dataa(Mux80),
	.datab(Mux16),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~29_cout ),
	.combout(),
	.cout(\LessThan1~31_cout ));
// synopsys translate_off
defparam \LessThan1~31 .lut_mask = 16'h004D;
defparam \LessThan1~31 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N0
cycloneive_lcell_comb \LessThan1~33 (
// Equation(s):
// \LessThan1~33_cout  = CARRY((\Mux79~0_combout  & ((!\LessThan1~31_cout ) # (!\Mux15~1_combout ))) # (!\Mux79~0_combout  & (!\Mux15~1_combout  & !\LessThan1~31_cout )))

	.dataa(Mux79),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~31_cout ),
	.combout(),
	.cout(\LessThan1~33_cout ));
// synopsys translate_off
defparam \LessThan1~33 .lut_mask = 16'h002B;
defparam \LessThan1~33 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N2
cycloneive_lcell_comb \LessThan1~35 (
// Equation(s):
// \LessThan1~35_cout  = CARRY((\Mux78~0_combout  & (\Mux14~1_combout  & !\LessThan1~33_cout )) # (!\Mux78~0_combout  & ((\Mux14~1_combout ) # (!\LessThan1~33_cout ))))

	.dataa(Mux78),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~33_cout ),
	.combout(),
	.cout(\LessThan1~35_cout ));
// synopsys translate_off
defparam \LessThan1~35 .lut_mask = 16'h004D;
defparam \LessThan1~35 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N4
cycloneive_lcell_comb \LessThan1~37 (
// Equation(s):
// \LessThan1~37_cout  = CARRY((\Mux13~1_combout  & (\Mux77~0_combout  & !\LessThan1~35_cout )) # (!\Mux13~1_combout  & ((\Mux77~0_combout ) # (!\LessThan1~35_cout ))))

	.dataa(Mux13),
	.datab(Mux77),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~35_cout ),
	.combout(),
	.cout(\LessThan1~37_cout ));
// synopsys translate_off
defparam \LessThan1~37 .lut_mask = 16'h004D;
defparam \LessThan1~37 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N6
cycloneive_lcell_comb \LessThan1~39 (
// Equation(s):
// \LessThan1~39_cout  = CARRY((\Mux76~0_combout  & (\Mux12~1_combout  & !\LessThan1~37_cout )) # (!\Mux76~0_combout  & ((\Mux12~1_combout ) # (!\LessThan1~37_cout ))))

	.dataa(Mux76),
	.datab(Mux12),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~37_cout ),
	.combout(),
	.cout(\LessThan1~39_cout ));
// synopsys translate_off
defparam \LessThan1~39 .lut_mask = 16'h004D;
defparam \LessThan1~39 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N8
cycloneive_lcell_comb \LessThan1~41 (
// Equation(s):
// \LessThan1~41_cout  = CARRY((\Mux11~1_combout  & (\Mux75~0_combout  & !\LessThan1~39_cout )) # (!\Mux11~1_combout  & ((\Mux75~0_combout ) # (!\LessThan1~39_cout ))))

	.dataa(Mux11),
	.datab(Mux75),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~39_cout ),
	.combout(),
	.cout(\LessThan1~41_cout ));
// synopsys translate_off
defparam \LessThan1~41 .lut_mask = 16'h004D;
defparam \LessThan1~41 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N10
cycloneive_lcell_comb \LessThan1~43 (
// Equation(s):
// \LessThan1~43_cout  = CARRY((\Mux10~1_combout  & ((!\LessThan1~41_cout ) # (!\Mux74~0_combout ))) # (!\Mux10~1_combout  & (!\Mux74~0_combout  & !\LessThan1~41_cout )))

	.dataa(Mux10),
	.datab(Mux74),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~41_cout ),
	.combout(),
	.cout(\LessThan1~43_cout ));
// synopsys translate_off
defparam \LessThan1~43 .lut_mask = 16'h002B;
defparam \LessThan1~43 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N12
cycloneive_lcell_comb \LessThan1~45 (
// Equation(s):
// \LessThan1~45_cout  = CARRY((\Mux9~1_combout  & (\Mux73~0_combout  & !\LessThan1~43_cout )) # (!\Mux9~1_combout  & ((\Mux73~0_combout ) # (!\LessThan1~43_cout ))))

	.dataa(Mux9),
	.datab(Mux73),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~43_cout ),
	.combout(),
	.cout(\LessThan1~45_cout ));
// synopsys translate_off
defparam \LessThan1~45 .lut_mask = 16'h004D;
defparam \LessThan1~45 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N14
cycloneive_lcell_comb \LessThan1~47 (
// Equation(s):
// \LessThan1~47_cout  = CARRY((\Mux8~1_combout  & ((!\LessThan1~45_cout ) # (!\Mux72~0_combout ))) # (!\Mux8~1_combout  & (!\Mux72~0_combout  & !\LessThan1~45_cout )))

	.dataa(Mux8),
	.datab(Mux72),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~45_cout ),
	.combout(),
	.cout(\LessThan1~47_cout ));
// synopsys translate_off
defparam \LessThan1~47 .lut_mask = 16'h002B;
defparam \LessThan1~47 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N16
cycloneive_lcell_comb \LessThan1~49 (
// Equation(s):
// \LessThan1~49_cout  = CARRY((\Mux7~1_combout  & (\Mux71~0_combout  & !\LessThan1~47_cout )) # (!\Mux7~1_combout  & ((\Mux71~0_combout ) # (!\LessThan1~47_cout ))))

	.dataa(Mux7),
	.datab(Mux71),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~47_cout ),
	.combout(),
	.cout(\LessThan1~49_cout ));
// synopsys translate_off
defparam \LessThan1~49 .lut_mask = 16'h004D;
defparam \LessThan1~49 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N18
cycloneive_lcell_comb \LessThan1~51 (
// Equation(s):
// \LessThan1~51_cout  = CARRY((\Mux6~1_combout  & ((!\LessThan1~49_cout ) # (!\Mux70~0_combout ))) # (!\Mux6~1_combout  & (!\Mux70~0_combout  & !\LessThan1~49_cout )))

	.dataa(Mux6),
	.datab(Mux70),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~49_cout ),
	.combout(),
	.cout(\LessThan1~51_cout ));
// synopsys translate_off
defparam \LessThan1~51 .lut_mask = 16'h002B;
defparam \LessThan1~51 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N20
cycloneive_lcell_comb \LessThan1~53 (
// Equation(s):
// \LessThan1~53_cout  = CARRY((\Mux5~1_combout  & (\Mux69~0_combout  & !\LessThan1~51_cout )) # (!\Mux5~1_combout  & ((\Mux69~0_combout ) # (!\LessThan1~51_cout ))))

	.dataa(Mux5),
	.datab(Mux69),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~51_cout ),
	.combout(),
	.cout(\LessThan1~53_cout ));
// synopsys translate_off
defparam \LessThan1~53 .lut_mask = 16'h004D;
defparam \LessThan1~53 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N22
cycloneive_lcell_comb \LessThan1~55 (
// Equation(s):
// \LessThan1~55_cout  = CARRY((\Mux68~0_combout  & (\Mux4~1_combout  & !\LessThan1~53_cout )) # (!\Mux68~0_combout  & ((\Mux4~1_combout ) # (!\LessThan1~53_cout ))))

	.dataa(Mux68),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~53_cout ),
	.combout(),
	.cout(\LessThan1~55_cout ));
// synopsys translate_off
defparam \LessThan1~55 .lut_mask = 16'h004D;
defparam \LessThan1~55 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N24
cycloneive_lcell_comb \LessThan1~57 (
// Equation(s):
// \LessThan1~57_cout  = CARRY((\Mux67~0_combout  & ((!\LessThan1~55_cout ) # (!\Mux3~1_combout ))) # (!\Mux67~0_combout  & (!\Mux3~1_combout  & !\LessThan1~55_cout )))

	.dataa(Mux67),
	.datab(Mux3),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~55_cout ),
	.combout(),
	.cout(\LessThan1~57_cout ));
// synopsys translate_off
defparam \LessThan1~57 .lut_mask = 16'h002B;
defparam \LessThan1~57 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N26
cycloneive_lcell_comb \LessThan1~59 (
// Equation(s):
// \LessThan1~59_cout  = CARRY((\Mux2~1_combout  & ((!\LessThan1~57_cout ) # (!\Mux66~0_combout ))) # (!\Mux2~1_combout  & (!\Mux66~0_combout  & !\LessThan1~57_cout )))

	.dataa(Mux2),
	.datab(Mux66),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~57_cout ),
	.combout(),
	.cout(\LessThan1~59_cout ));
// synopsys translate_off
defparam \LessThan1~59 .lut_mask = 16'h002B;
defparam \LessThan1~59 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N28
cycloneive_lcell_comb \LessThan1~61 (
// Equation(s):
// \LessThan1~61_cout  = CARRY((\Mux65~0_combout  & ((!\LessThan1~59_cout ) # (!\Mux1~1_combout ))) # (!\Mux65~0_combout  & (!\Mux1~1_combout  & !\LessThan1~59_cout )))

	.dataa(Mux65),
	.datab(Mux1),
	.datac(gnd),
	.datad(vcc),
	.cin(\LessThan1~59_cout ),
	.combout(),
	.cout(\LessThan1~61_cout ));
// synopsys translate_off
defparam \LessThan1~61 .lut_mask = 16'h002B;
defparam \LessThan1~61 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X53_Y23_N30
cycloneive_lcell_comb \LessThan1~62 (
// Equation(s):
// \LessThan1~62_combout  = (\Mux0~1_combout  & (\LessThan1~61_cout  & \Mux64~0_combout )) # (!\Mux0~1_combout  & ((\LessThan1~61_cout ) # (\Mux64~0_combout )))

	.dataa(gnd),
	.datab(Mux0),
	.datac(gnd),
	.datad(Mux64),
	.cin(\LessThan1~61_cout ),
	.combout(\LessThan1~62_combout ),
	.cout());
// synopsys translate_off
defparam \LessThan1~62 .lut_mask = 16'hF330;
defparam \LessThan1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N24
cycloneive_lcell_comb \aluif.portOut[0]~23 (
// Equation(s):
// \aluif.portOut[0]~23_combout  = (\prif.ALUOP_ex [2] & ((\prif.ALUOP_ex [0] & (\LessThan0~62_combout )) # (!\prif.ALUOP_ex [0] & ((\LessThan1~62_combout )))))

	.dataa(\LessThan0~62_combout ),
	.datab(prifALUOP_ex_0),
	.datac(\LessThan1~62_combout ),
	.datad(prifALUOP_ex_2),
	.cin(gnd),
	.combout(\aluif.portOut[0]~23_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[0]~23 .lut_mask = 16'hB800;
defparam \aluif.portOut[0]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N22
cycloneive_lcell_comb \portOut~4 (
// Equation(s):
// \portOut~4_combout  = (\Mux28~1_combout ) # (\Mux92~2_combout )

	.dataa(Mux28),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux92),
	.cin(gnd),
	.combout(\portOut~4_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~4 .lut_mask = 16'hFFAA;
defparam \portOut~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N20
cycloneive_lcell_comb \aluif.portOut[5]~25 (
// Equation(s):
// \aluif.portOut[5]~25_combout  = (\prif.ALUOP_ex [3] & \prif.ALUOP_ex [0])

	.dataa(gnd),
	.datab(gnd),
	.datac(prifALUOP_ex_3),
	.datad(prifALUOP_ex_0),
	.cin(gnd),
	.combout(\aluif.portOut[5]~25_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~25 .lut_mask = 16'hF000;
defparam \aluif.portOut[5]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N4
cycloneive_lcell_comb \aluif.portOut[2]~29 (
// Equation(s):
// \aluif.portOut[2]~29_combout  = (\prif.ALUOP_ex [3] & (!\prif.ALUOP_ex [1] & (!\prif.ALUOP_ex [0] & !\prif.ALUOP_ex [2])))

	.dataa(prifALUOP_ex_3),
	.datab(prifALUOP_ex_1),
	.datac(prifALUOP_ex_0),
	.datad(prifALUOP_ex_2),
	.cin(gnd),
	.combout(\aluif.portOut[2]~29_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~29 .lut_mask = 16'h0002;
defparam \aluif.portOut[2]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N4
cycloneive_lcell_comb \Add0~4 (
// Equation(s):
// \Add0~4_combout  = ((\Mux29~1_combout  $ (\Mux93~2_combout  $ (!\Add0~3 )))) # (GND)
// \Add0~5  = CARRY((\Mux29~1_combout  & ((\Mux93~2_combout ) # (!\Add0~3 ))) # (!\Mux29~1_combout  & (\Mux93~2_combout  & !\Add0~3 )))

	.dataa(Mux29),
	.datab(Mux931),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~3 ),
	.combout(\Add0~4_combout ),
	.cout(\Add0~5 ));
// synopsys translate_off
defparam \Add0~4 .lut_mask = 16'h698E;
defparam \Add0~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N6
cycloneive_lcell_comb \Add0~6 (
// Equation(s):
// \Add0~6_combout  = (\Mux28~1_combout  & ((\Mux92~2_combout  & (\Add0~5  & VCC)) # (!\Mux92~2_combout  & (!\Add0~5 )))) # (!\Mux28~1_combout  & ((\Mux92~2_combout  & (!\Add0~5 )) # (!\Mux92~2_combout  & ((\Add0~5 ) # (GND)))))
// \Add0~7  = CARRY((\Mux28~1_combout  & (!\Mux92~2_combout  & !\Add0~5 )) # (!\Mux28~1_combout  & ((!\Add0~5 ) # (!\Mux92~2_combout ))))

	.dataa(Mux28),
	.datab(Mux92),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~5 ),
	.combout(\Add0~6_combout ),
	.cout(\Add0~7 ));
// synopsys translate_off
defparam \Add0~6 .lut_mask = 16'h9617;
defparam \Add0~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N0
cycloneive_lcell_comb \portOut~2 (
// Equation(s):
// \portOut~2_combout  = \Mux28~1_combout  $ (\Mux92~2_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux28),
	.datad(Mux92),
	.cin(gnd),
	.combout(\portOut~2_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~2 .lut_mask = 16'h0FF0;
defparam \portOut~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N18
cycloneive_lcell_comb \aluif.portOut[15]~26 (
// Equation(s):
// \aluif.portOut[15]~26_combout  = (\prif.ALUOP_ex [1] & (((!\ShiftLeft0~15_combout  & !\Mux91~2_combout )) # (!\prif.ALUOP_ex [2])))

	.dataa(prifALUOP_ex_2),
	.datab(prifALUOP_ex_1),
	.datac(\ShiftLeft0~15_combout ),
	.datad(Mux91),
	.cin(gnd),
	.combout(\aluif.portOut[15]~26_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~26 .lut_mask = 16'h444C;
defparam \aluif.portOut[15]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y22_N2
cycloneive_lcell_comb \portOut~3 (
// Equation(s):
// \portOut~3_combout  = (\Mux92~2_combout  & \Mux28~1_combout )

	.dataa(gnd),
	.datab(Mux92),
	.datac(gnd),
	.datad(Mux28),
	.cin(gnd),
	.combout(\portOut~3_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~3 .lut_mask = 16'hCC00;
defparam \portOut~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y22_N12
cycloneive_lcell_comb \aluif.portOut[3]~27 (
// Equation(s):
// \aluif.portOut[3]~27_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & (\ShiftLeft0~19_combout )) # (!\prif.ALUOP_ex [2] & ((\portOut~3_combout ))))) # (!\aluif.portOut[15]~26_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\ShiftLeft0~19_combout ),
	.datab(\aluif.portOut[15]~26_combout ),
	.datac(prifALUOP_ex_2),
	.datad(\portOut~3_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[3]~27_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[3]~27 .lut_mask = 16'h8F83;
defparam \aluif.portOut[3]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y22_N30
cycloneive_lcell_comb \aluif.portOut[3]~28 (
// Equation(s):
// \aluif.portOut[3]~28_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[3]~27_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[3]~27_combout  & ((\portOut~2_combout ))) # (!\aluif.portOut[3]~27_combout  & (\Add0~6_combout ))))

	.dataa(\Add0~6_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\portOut~2_combout ),
	.datad(\aluif.portOut[3]~27_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[3]~28_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[3]~28 .lut_mask = 16'hFC22;
defparam \aluif.portOut[3]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N12
cycloneive_lcell_comb \aluif.portOut[2]~32 (
// Equation(s):
// \aluif.portOut[2]~32_combout  = (!\prif.ALUOP_ex [2] & !\prif.ALUOP_ex [1])

	.dataa(gnd),
	.datab(prifALUOP_ex_2),
	.datac(gnd),
	.datad(prifALUOP_ex_1),
	.cin(gnd),
	.combout(\aluif.portOut[2]~32_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~32 .lut_mask = 16'h0033;
defparam \aluif.portOut[2]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N4
cycloneive_lcell_comb \Add1~4 (
// Equation(s):
// \Add1~4_combout  = ((\Mux29~1_combout  $ (\Mux93~2_combout  $ (\Add1~3 )))) # (GND)
// \Add1~5  = CARRY((\Mux29~1_combout  & ((!\Add1~3 ) # (!\Mux93~2_combout ))) # (!\Mux29~1_combout  & (!\Mux93~2_combout  & !\Add1~3 )))

	.dataa(Mux29),
	.datab(Mux931),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'h962B;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N6
cycloneive_lcell_comb \Add1~6 (
// Equation(s):
// \Add1~6_combout  = (\Mux28~1_combout  & ((\Mux92~2_combout  & (!\Add1~5 )) # (!\Mux92~2_combout  & (\Add1~5  & VCC)))) # (!\Mux28~1_combout  & ((\Mux92~2_combout  & ((\Add1~5 ) # (GND))) # (!\Mux92~2_combout  & (!\Add1~5 ))))
// \Add1~7  = CARRY((\Mux28~1_combout  & (\Mux92~2_combout  & !\Add1~5 )) # (!\Mux28~1_combout  & ((\Mux92~2_combout ) # (!\Add1~5 ))))

	.dataa(Mux28),
	.datab(Mux92),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h694D;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N16
cycloneive_lcell_comb \aluif.portOut[2]~34 (
// Equation(s):
// \aluif.portOut[2]~34_combout  = ((\prif.ALUOP_ex [2] & \Mux91~2_combout )) # (!\prif.ALUOP_ex [1])

	.dataa(prifALUOP_ex_2),
	.datab(prifALUOP_ex_1),
	.datac(gnd),
	.datad(Mux91),
	.cin(gnd),
	.combout(\aluif.portOut[2]~34_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~34 .lut_mask = 16'hBB33;
defparam \aluif.portOut[2]~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N20
cycloneive_lcell_comb \aluif.portOut[2]~35 (
// Equation(s):
// \aluif.portOut[2]~35_combout  = (\Mux92~2_combout ) # ((\Mux94~1_combout  & !\Mux93~2_combout ))

	.dataa(gnd),
	.datab(Mux94),
	.datac(Mux931),
	.datad(Mux92),
	.cin(gnd),
	.combout(\aluif.portOut[2]~35_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~35 .lut_mask = 16'hFF0C;
defparam \aluif.portOut[2]~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N16
cycloneive_lcell_comb \ShiftRight0~10 (
// Equation(s):
// \ShiftRight0~10_combout  = (\Mux95~1_combout  & ((\Mux25~1_combout ))) # (!\Mux95~1_combout  & (\Mux26~1_combout ))

	.dataa(gnd),
	.datab(Mux26),
	.datac(Mux25),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~10_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~10 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N16
cycloneive_lcell_comb \ShiftRight0~61 (
// Equation(s):
// \ShiftRight0~61_combout  = (!\Mux93~2_combout  & !\Mux92~2_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux931),
	.datad(Mux92),
	.cin(gnd),
	.combout(\ShiftRight0~61_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~61 .lut_mask = 16'h000F;
defparam \ShiftRight0~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N14
cycloneive_lcell_comb \ShiftRight0~17 (
// Equation(s):
// \ShiftRight0~17_combout  = (\Mux95~1_combout  & (\Mux21~1_combout )) # (!\Mux95~1_combout  & ((\Mux22~1_combout )))

	.dataa(Mux21),
	.datab(Mux22),
	.datac(gnd),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~17 .lut_mask = 16'hAACC;
defparam \ShiftRight0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N16
cycloneive_lcell_comb \ShiftRight0~9 (
// Equation(s):
// \ShiftRight0~9_combout  = (\Mux95~1_combout  & ((\Mux23~1_combout ))) # (!\Mux95~1_combout  & (\Mux24~1_combout ))

	.dataa(Mux24),
	.datab(gnd),
	.datac(Mux23),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~9_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~9 .lut_mask = 16'hF0AA;
defparam \ShiftRight0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N26
cycloneive_lcell_comb \ShiftRight0~72 (
// Equation(s):
// \ShiftRight0~72_combout  = (\Mux94~1_combout  & (\ShiftRight0~17_combout )) # (!\Mux94~1_combout  & ((\ShiftRight0~9_combout )))

	.dataa(Mux94),
	.datab(\ShiftRight0~17_combout ),
	.datac(\ShiftRight0~9_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~72 .lut_mask = 16'hD8D8;
defparam \ShiftRight0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N12
cycloneive_lcell_comb \ShiftRight0~7 (
// Equation(s):
// \ShiftRight0~7_combout  = (\Mux95~1_combout  & ((\Mux27~1_combout ))) # (!\Mux95~1_combout  & (\Mux28~1_combout ))

	.dataa(gnd),
	.datab(Mux28),
	.datac(Mux27),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~7_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~7 .lut_mask = 16'hF0CC;
defparam \ShiftRight0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N20
cycloneive_lcell_comb \aluif.portOut[3]~36 (
// Equation(s):
// \aluif.portOut[3]~36_combout  = (\aluif.portOut[2]~35_combout  & (!\ShiftRight0~61_combout )) # (!\aluif.portOut[2]~35_combout  & ((\ShiftRight0~61_combout  & ((\ShiftRight0~7_combout ))) # (!\ShiftRight0~61_combout  & (\ShiftRight0~72_combout ))))

	.dataa(\aluif.portOut[2]~35_combout ),
	.datab(\ShiftRight0~61_combout ),
	.datac(\ShiftRight0~72_combout ),
	.datad(\ShiftRight0~7_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[3]~36_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[3]~36 .lut_mask = 16'h7632;
defparam \aluif.portOut[3]~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N14
cycloneive_lcell_comb \aluif.portOut[3]~37 (
// Equation(s):
// \aluif.portOut[3]~37_combout  = (\aluif.portOut[2]~35_combout  & ((\aluif.portOut[3]~36_combout  & (\ShiftRight0~76_combout )) # (!\aluif.portOut[3]~36_combout  & ((\ShiftRight0~10_combout ))))) # (!\aluif.portOut[2]~35_combout  & 
// (((\aluif.portOut[3]~36_combout ))))

	.dataa(\ShiftRight0~76_combout ),
	.datab(\aluif.portOut[2]~35_combout ),
	.datac(\ShiftRight0~10_combout ),
	.datad(\aluif.portOut[3]~36_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[3]~37_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[3]~37 .lut_mask = 16'hBBC0;
defparam \aluif.portOut[3]~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N20
cycloneive_lcell_comb \ShiftRight0~62 (
// Equation(s):
// \ShiftRight0~62_combout  = (\Mux0~1_combout  & (!\Mux95~1_combout  & !\Mux94~1_combout ))

	.dataa(Mux0),
	.datab(gnd),
	.datac(Mux95),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftRight0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~62 .lut_mask = 16'h000A;
defparam \ShiftRight0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N26
cycloneive_lcell_comb \ShiftRight0~63 (
// Equation(s):
// \ShiftRight0~63_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux1~1_combout ))) # (!\Mux95~1_combout  & (\Mux2~1_combout ))))

	.dataa(Mux2),
	.datab(Mux94),
	.datac(Mux95),
	.datad(Mux1),
	.cin(gnd),
	.combout(\ShiftRight0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~63 .lut_mask = 16'hC808;
defparam \ShiftRight0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N4
cycloneive_lcell_comb \ShiftRight0~65 (
// Equation(s):
// \ShiftRight0~65_combout  = (\Mux93~2_combout  & (((\ShiftRight0~62_combout )))) # (!\Mux93~2_combout  & ((\ShiftRight0~64_combout ) # ((\ShiftRight0~63_combout ))))

	.dataa(\ShiftRight0~64_combout ),
	.datab(\ShiftRight0~62_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~63_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~65 .lut_mask = 16'hCFCA;
defparam \ShiftRight0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N8
cycloneive_lcell_comb \ShiftRight0~66 (
// Equation(s):
// \ShiftRight0~66_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux5~1_combout )) # (!\Mux95~1_combout  & ((\Mux6~1_combout ))))) # (!\Mux94~1_combout  & (((\Mux95~1_combout ))))

	.dataa(Mux94),
	.datab(Mux5),
	.datac(Mux95),
	.datad(Mux6),
	.cin(gnd),
	.combout(\ShiftRight0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~66 .lut_mask = 16'hDAD0;
defparam \ShiftRight0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N14
cycloneive_lcell_comb \ShiftRight0~67 (
// Equation(s):
// \ShiftRight0~67_combout  = (\ShiftRight0~66_combout  & ((\Mux7~1_combout ) # ((\Mux94~1_combout )))) # (!\ShiftRight0~66_combout  & (((\Mux8~1_combout  & !\Mux94~1_combout ))))

	.dataa(Mux7),
	.datab(Mux8),
	.datac(\ShiftRight0~66_combout ),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftRight0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~67 .lut_mask = 16'hF0AC;
defparam \ShiftRight0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N10
cycloneive_lcell_comb \ShiftRight0~70 (
// Equation(s):
// \ShiftRight0~70_combout  = (\Mux93~2_combout  & ((\ShiftRight0~67_combout ))) # (!\Mux93~2_combout  & (\ShiftRight0~69_combout ))

	.dataa(\ShiftRight0~69_combout ),
	.datab(gnd),
	.datac(Mux931),
	.datad(\ShiftRight0~67_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~70 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N8
cycloneive_lcell_comb \ShiftRight0~71 (
// Equation(s):
// \ShiftRight0~71_combout  = (\Mux92~2_combout  & (\ShiftRight0~65_combout )) # (!\Mux92~2_combout  & ((\ShiftRight0~70_combout )))

	.dataa(gnd),
	.datab(Mux92),
	.datac(\ShiftRight0~65_combout ),
	.datad(\ShiftRight0~70_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~71 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N0
cycloneive_lcell_comb \aluif.portOut[3]~38 (
// Equation(s):
// \aluif.portOut[3]~38_combout  = (\aluif.portOut[1]~13_combout  & ((\aluif.portOut[2]~34_combout  & ((\ShiftRight0~71_combout ))) # (!\aluif.portOut[2]~34_combout  & (\aluif.portOut[3]~37_combout )))) # (!\aluif.portOut[1]~13_combout  & 
// (\aluif.portOut[2]~34_combout ))

	.dataa(\aluif.portOut[1]~13_combout ),
	.datab(\aluif.portOut[2]~34_combout ),
	.datac(\aluif.portOut[3]~37_combout ),
	.datad(\ShiftRight0~71_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[3]~38_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[3]~38 .lut_mask = 16'hEC64;
defparam \aluif.portOut[3]~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N24
cycloneive_lcell_comb \ShiftRight0~90 (
// Equation(s):
// \ShiftRight0~90_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux14~1_combout )) # (!\Mux95~1_combout  & ((\Mux15~1_combout )))))

	.dataa(Mux94),
	.datab(Mux95),
	.datac(Mux14),
	.datad(Mux15),
	.cin(gnd),
	.combout(\ShiftRight0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~90 .lut_mask = 16'hA280;
defparam \ShiftRight0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N16
cycloneive_lcell_comb \ShiftRight0~88 (
// Equation(s):
// \ShiftRight0~88_combout  = (\Mux94~1_combout  & (\ShiftRight0~54_combout )) # (!\Mux94~1_combout  & ((\ShiftRight0~56_combout )))

	.dataa(gnd),
	.datab(\ShiftRight0~54_combout ),
	.datac(Mux94),
	.datad(\ShiftRight0~56_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~88 .lut_mask = 16'hCFC0;
defparam \ShiftRight0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N14
cycloneive_lcell_comb \ShiftRight0~91 (
// Equation(s):
// \ShiftRight0~91_combout  = (\Mux93~2_combout  & ((\ShiftRight0~89_combout ) # ((\ShiftRight0~90_combout )))) # (!\Mux93~2_combout  & (((\ShiftRight0~88_combout ))))

	.dataa(\ShiftRight0~89_combout ),
	.datab(\ShiftRight0~90_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~88_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~91 .lut_mask = 16'hEFE0;
defparam \ShiftRight0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N2
cycloneive_lcell_comb \ShiftRight0~87 (
// Equation(s):
// \ShiftRight0~87_combout  = (\Mux94~1_combout  & ((\ShiftRight0~57_combout ))) # (!\Mux94~1_combout  & (\ShiftRight0~49_combout ))

	.dataa(\ShiftRight0~49_combout ),
	.datab(gnd),
	.datac(Mux94),
	.datad(\ShiftRight0~57_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~87 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N28
cycloneive_lcell_comb \aluif.portOut[2]~44 (
// Equation(s):
// \aluif.portOut[2]~44_combout  = (\aluif.portOut[2]~35_combout  & (((!\ShiftRight0~61_combout )))) # (!\aluif.portOut[2]~35_combout  & ((\ShiftRight0~61_combout  & ((\ShiftRight0~47_combout ))) # (!\ShiftRight0~61_combout  & (\ShiftRight0~87_combout ))))

	.dataa(\aluif.portOut[2]~35_combout ),
	.datab(\ShiftRight0~87_combout ),
	.datac(\ShiftRight0~61_combout ),
	.datad(\ShiftRight0~47_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[2]~44_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~44 .lut_mask = 16'h5E0E;
defparam \aluif.portOut[2]~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N12
cycloneive_lcell_comb \aluif.portOut[2]~45 (
// Equation(s):
// \aluif.portOut[2]~45_combout  = (\aluif.portOut[2]~35_combout  & ((\aluif.portOut[2]~44_combout  & ((\ShiftRight0~91_combout ))) # (!\aluif.portOut[2]~44_combout  & (\ShiftRight0~50_combout )))) # (!\aluif.portOut[2]~35_combout  & 
// (((\aluif.portOut[2]~44_combout ))))

	.dataa(\aluif.portOut[2]~35_combout ),
	.datab(\ShiftRight0~50_combout ),
	.datac(\ShiftRight0~91_combout ),
	.datad(\aluif.portOut[2]~44_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[2]~45_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~45 .lut_mask = 16'hF588;
defparam \aluif.portOut[2]~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N24
cycloneive_lcell_comb \portOut~7 (
// Equation(s):
// \portOut~7_combout  = (\Mux93~2_combout ) # (\Mux29~1_combout )

	.dataa(gnd),
	.datab(Mux931),
	.datac(Mux29),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~7_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~7 .lut_mask = 16'hFCFC;
defparam \portOut~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N20
cycloneive_lcell_comb \aluif.portOut[2]~46 (
// Equation(s):
// \aluif.portOut[2]~46_combout  = (\aluif.portOut[1]~13_combout  & (!\aluif.portOut[2]~34_combout  & (\aluif.portOut[2]~45_combout ))) # (!\aluif.portOut[1]~13_combout  & ((\aluif.portOut[2]~34_combout ) # ((\portOut~7_combout ))))

	.dataa(\aluif.portOut[1]~13_combout ),
	.datab(\aluif.portOut[2]~34_combout ),
	.datac(\aluif.portOut[2]~45_combout ),
	.datad(\portOut~7_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[2]~46_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~46 .lut_mask = 16'h7564;
defparam \aluif.portOut[2]~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N24
cycloneive_lcell_comb \ShiftRight0~77 (
// Equation(s):
// \ShiftRight0~77_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux0~1_combout ))) # (!\Mux95~1_combout  & (\Mux1~1_combout ))))

	.dataa(Mux1),
	.datab(Mux95),
	.datac(Mux0),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftRight0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~77 .lut_mask = 16'h00E2;
defparam \ShiftRight0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N30
cycloneive_lcell_comb \ShiftRight0~80 (
// Equation(s):
// \ShiftRight0~80_combout  = (\Mux92~2_combout  & ((\Mux93~2_combout  & ((\ShiftRight0~77_combout ))) # (!\Mux93~2_combout  & (\ShiftRight0~79_combout ))))

	.dataa(\ShiftRight0~79_combout ),
	.datab(Mux92),
	.datac(Mux931),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~80 .lut_mask = 16'hC808;
defparam \ShiftRight0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N8
cycloneive_lcell_comb \ShiftRight0~81 (
// Equation(s):
// \ShiftRight0~81_combout  = (\Mux95~1_combout  & (((\Mux6~1_combout )) # (!\Mux94~1_combout ))) # (!\Mux95~1_combout  & (\Mux94~1_combout  & ((\Mux7~1_combout ))))

	.dataa(Mux95),
	.datab(Mux94),
	.datac(Mux6),
	.datad(Mux7),
	.cin(gnd),
	.combout(\ShiftRight0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~81 .lut_mask = 16'hE6A2;
defparam \ShiftRight0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N18
cycloneive_lcell_comb \ShiftRight0~82 (
// Equation(s):
// \ShiftRight0~82_combout  = (\Mux94~1_combout  & (((\ShiftRight0~81_combout )))) # (!\Mux94~1_combout  & ((\ShiftRight0~81_combout  & ((\Mux8~1_combout ))) # (!\ShiftRight0~81_combout  & (\Mux9~1_combout ))))

	.dataa(Mux9),
	.datab(Mux94),
	.datac(\ShiftRight0~81_combout ),
	.datad(Mux8),
	.cin(gnd),
	.combout(\ShiftRight0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~82 .lut_mask = 16'hF2C2;
defparam \ShiftRight0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N28
cycloneive_lcell_comb \ShiftRight0~85 (
// Equation(s):
// \ShiftRight0~85_combout  = (\Mux93~2_combout  & ((\ShiftRight0~82_combout ))) # (!\Mux93~2_combout  & (\ShiftRight0~84_combout ))

	.dataa(\ShiftRight0~84_combout ),
	.datab(gnd),
	.datac(Mux931),
	.datad(\ShiftRight0~82_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~85 .lut_mask = 16'hFA0A;
defparam \ShiftRight0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N26
cycloneive_lcell_comb \ShiftRight0~86 (
// Equation(s):
// \ShiftRight0~86_combout  = (\ShiftRight0~80_combout ) # ((!\Mux92~2_combout  & \ShiftRight0~85_combout ))

	.dataa(gnd),
	.datab(Mux92),
	.datac(\ShiftRight0~80_combout ),
	.datad(\ShiftRight0~85_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~86 .lut_mask = 16'hF3F0;
defparam \ShiftRight0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N18
cycloneive_lcell_comb \aluif.portOut[2]~47 (
// Equation(s):
// \aluif.portOut[2]~47_combout  = (\aluif.portOut[2]~34_combout  & ((\aluif.portOut[2]~46_combout  & (\Add1~4_combout )) # (!\aluif.portOut[2]~46_combout  & ((\ShiftRight0~86_combout ))))) # (!\aluif.portOut[2]~34_combout  & (((\aluif.portOut[2]~46_combout 
// ))))

	.dataa(\Add1~4_combout ),
	.datab(\aluif.portOut[2]~34_combout ),
	.datac(\aluif.portOut[2]~46_combout ),
	.datad(\ShiftRight0~86_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[2]~47_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~47 .lut_mask = 16'hBCB0;
defparam \aluif.portOut[2]~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N20
cycloneive_lcell_comb \ShiftLeft0~20 (
// Equation(s):
// \ShiftLeft0~20_combout  = (!\Mux95~1_combout  & ((\Mux94~1_combout  & ((\Mux31~1_combout ))) # (!\Mux94~1_combout  & (\Mux29~1_combout ))))

	.dataa(Mux29),
	.datab(Mux95),
	.datac(Mux31),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftLeft0~20_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~20 .lut_mask = 16'h3022;
defparam \ShiftLeft0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N2
cycloneive_lcell_comb \ShiftLeft0~21 (
// Equation(s):
// \ShiftLeft0~21_combout  = (\ShiftLeft0~20_combout ) # ((!\Mux94~1_combout  & (\Mux30~1_combout  & \Mux95~1_combout )))

	.dataa(Mux94),
	.datab(Mux30),
	.datac(Mux95),
	.datad(\ShiftLeft0~20_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~21_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~21 .lut_mask = 16'hFF40;
defparam \ShiftLeft0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N30
cycloneive_lcell_comb \ShiftLeft0~109 (
// Equation(s):
// \ShiftLeft0~109_combout  = (!\Mux93~2_combout  & (!\Mux92~2_combout  & \ShiftLeft0~21_combout ))

	.dataa(Mux931),
	.datab(gnd),
	.datac(Mux92),
	.datad(\ShiftLeft0~21_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~109_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~109 .lut_mask = 16'h0500;
defparam \ShiftLeft0~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N16
cycloneive_lcell_comb \aluif.portOut[2]~41 (
// Equation(s):
// \aluif.portOut[2]~41_combout  = (\prif.ALUOP_ex [2] & (((\ShiftLeft0~109_combout  & \aluif.portOut[15]~26_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~6_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(\portOut~6_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\ShiftLeft0~109_combout ),
	.datad(\aluif.portOut[15]~26_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[2]~41_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~41 .lut_mask = 16'hE233;
defparam \aluif.portOut[2]~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N26
cycloneive_lcell_comb \aluif.portOut[2]~42 (
// Equation(s):
// \aluif.portOut[2]~42_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[2]~41_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[2]~41_combout  & (\portOut~5_combout )) # (!\aluif.portOut[2]~41_combout  & ((\Add0~4_combout )))))

	.dataa(\portOut~5_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\Add0~4_combout ),
	.datad(\aluif.portOut[2]~41_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[2]~42_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~42 .lut_mask = 16'hEE30;
defparam \aluif.portOut[2]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N2
cycloneive_lcell_comb \aluif.portOut[2]~43 (
// Equation(s):
// \aluif.portOut[2]~43_combout  = (\aluif.portOut[2]~42_combout  & ((\aluif.portOut[5]~25_combout ) # ((!\portOut~7_combout  & \aluif.portOut[2]~29_combout )))) # (!\aluif.portOut[2]~42_combout  & (!\portOut~7_combout  & (\aluif.portOut[2]~29_combout )))

	.dataa(\aluif.portOut[2]~42_combout ),
	.datab(\portOut~7_combout ),
	.datac(\aluif.portOut[2]~29_combout ),
	.datad(\aluif.portOut[5]~25_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[2]~43_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[2]~43 .lut_mask = 16'hBA30;
defparam \aluif.portOut[2]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N8
cycloneive_lcell_comb \Add1~8 (
// Equation(s):
// \Add1~8_combout  = ((\Mux91~2_combout  $ (\Mux27~1_combout  $ (\Add1~7 )))) # (GND)
// \Add1~9  = CARRY((\Mux91~2_combout  & (\Mux27~1_combout  & !\Add1~7 )) # (!\Mux91~2_combout  & ((\Mux27~1_combout ) # (!\Add1~7 ))))

	.dataa(Mux91),
	.datab(Mux27),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'h964D;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N10
cycloneive_lcell_comb \Add1~10 (
// Equation(s):
// \Add1~10_combout  = (\Mux26~1_combout  & ((\Mux90~3_combout  & (!\Add1~9 )) # (!\Mux90~3_combout  & (\Add1~9  & VCC)))) # (!\Mux26~1_combout  & ((\Mux90~3_combout  & ((\Add1~9 ) # (GND))) # (!\Mux90~3_combout  & (!\Add1~9 ))))
// \Add1~11  = CARRY((\Mux26~1_combout  & (\Mux90~3_combout  & !\Add1~9 )) # (!\Mux26~1_combout  & ((\Mux90~3_combout ) # (!\Add1~9 ))))

	.dataa(Mux26),
	.datab(Mux90),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout(\Add1~11 ));
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h694D;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N12
cycloneive_lcell_comb \portOut~10 (
// Equation(s):
// \portOut~10_combout  = (\Mux90~3_combout ) # (\Mux26~1_combout )

	.dataa(gnd),
	.datab(Mux90),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\portOut~10_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~10 .lut_mask = 16'hFFCC;
defparam \portOut~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N10
cycloneive_lcell_comb \aluif.portOut[5]~55 (
// Equation(s):
// \aluif.portOut[5]~55_combout  = (\prif.ALUOP_ex [1] & ((!\prif.ALUOP_ex [2]) # (!\ShiftLeft0~15_combout )))

	.dataa(gnd),
	.datab(prifALUOP_ex_1),
	.datac(\ShiftLeft0~15_combout ),
	.datad(prifALUOP_ex_2),
	.cin(gnd),
	.combout(\aluif.portOut[5]~55_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~55 .lut_mask = 16'h0CCC;
defparam \aluif.portOut[5]~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N8
cycloneive_lcell_comb \aluif.portOut[5]~51 (
// Equation(s):
// \aluif.portOut[5]~51_combout  = (\Mux91~2_combout ) # (\Mux92~2_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux91),
	.datad(Mux92),
	.cin(gnd),
	.combout(\aluif.portOut[5]~51_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~51 .lut_mask = 16'hFFF0;
defparam \aluif.portOut[5]~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N8
cycloneive_lcell_comb \ShiftRight0~93 (
// Equation(s):
// \ShiftRight0~93_combout  = (\ShiftRight0~28_combout ) # (\ShiftRight0~29_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(\ShiftRight0~28_combout ),
	.datad(\ShiftRight0~29_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~93 .lut_mask = 16'hFFF0;
defparam \ShiftRight0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N12
cycloneive_lcell_comb \ShiftRight0~24 (
// Equation(s):
// \ShiftRight0~24_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux7~1_combout ))) # (!\Mux95~1_combout  & (\Mux8~1_combout ))))

	.dataa(Mux94),
	.datab(Mux95),
	.datac(Mux8),
	.datad(Mux7),
	.cin(gnd),
	.combout(\ShiftRight0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~24 .lut_mask = 16'hA820;
defparam \ShiftRight0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N14
cycloneive_lcell_comb \ShiftRight0~94 (
// Equation(s):
// \ShiftRight0~94_combout  = (\Mux93~2_combout  & (((\ShiftRight0~93_combout )))) # (!\Mux93~2_combout  & ((\ShiftRight0~23_combout ) # ((\ShiftRight0~24_combout ))))

	.dataa(Mux931),
	.datab(\ShiftRight0~23_combout ),
	.datac(\ShiftRight0~93_combout ),
	.datad(\ShiftRight0~24_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~94 .lut_mask = 16'hF5E4;
defparam \ShiftRight0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N10
cycloneive_lcell_comb \ShiftRight0~112 (
// Equation(s):
// \ShiftRight0~112_combout  = (\ShiftRight0~26_combout ) # ((!\Mux94~1_combout  & (!\Mux95~1_combout  & \Mux2~1_combout )))

	.dataa(Mux94),
	.datab(\ShiftRight0~26_combout ),
	.datac(Mux95),
	.datad(Mux2),
	.cin(gnd),
	.combout(\ShiftRight0~112_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~112 .lut_mask = 16'hCDCC;
defparam \ShiftRight0~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N12
cycloneive_lcell_comb \ShiftRight0~95 (
// Equation(s):
// \ShiftRight0~95_combout  = (\Mux92~2_combout  & (((!\Mux93~2_combout  & \ShiftRight0~112_combout )))) # (!\Mux92~2_combout  & (\ShiftRight0~94_combout ))

	.dataa(Mux92),
	.datab(\ShiftRight0~94_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~112_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~95_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~95 .lut_mask = 16'h4E44;
defparam \ShiftRight0~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N14
cycloneive_lcell_comb \ShiftRight0~14 (
// Equation(s):
// \ShiftRight0~14_combout  = (\Mux95~1_combout  & ((\Mux17~1_combout ))) # (!\Mux95~1_combout  & (\Mux18~1_combout ))

	.dataa(Mux18),
	.datab(Mux17),
	.datac(gnd),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~14_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~14 .lut_mask = 16'hCCAA;
defparam \ShiftRight0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N12
cycloneive_lcell_comb \ShiftRight0~13 (
// Equation(s):
// \ShiftRight0~13_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux15~1_combout )) # (!\Mux95~1_combout  & ((\Mux16~1_combout )))))

	.dataa(Mux15),
	.datab(Mux94),
	.datac(Mux16),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~13_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~13 .lut_mask = 16'h88C0;
defparam \ShiftRight0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N8
cycloneive_lcell_comb \ShiftRight0~15 (
// Equation(s):
// \ShiftRight0~15_combout  = (\ShiftRight0~13_combout ) # ((!\Mux94~1_combout  & \ShiftRight0~14_combout ))

	.dataa(gnd),
	.datab(Mux94),
	.datac(\ShiftRight0~14_combout ),
	.datad(\ShiftRight0~13_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~15_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~15 .lut_mask = 16'hFF30;
defparam \ShiftRight0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N20
cycloneive_lcell_comb \ShiftRight0~92 (
// Equation(s):
// \ShiftRight0~92_combout  = (\Mux93~2_combout  & ((\ShiftRight0~22_combout ))) # (!\Mux93~2_combout  & (\ShiftRight0~15_combout ))

	.dataa(gnd),
	.datab(Mux931),
	.datac(\ShiftRight0~15_combout ),
	.datad(\ShiftRight0~22_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~92 .lut_mask = 16'hFC30;
defparam \ShiftRight0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N2
cycloneive_lcell_comb \aluif.portOut[5]~54 (
// Equation(s):
// \aluif.portOut[5]~54_combout  = (\aluif.portOut[5]~53_combout  & (((\ShiftRight0~95_combout )) # (!\aluif.portOut[5]~51_combout ))) # (!\aluif.portOut[5]~53_combout  & (\aluif.portOut[5]~51_combout  & ((\ShiftRight0~92_combout ))))

	.dataa(\aluif.portOut[5]~53_combout ),
	.datab(\aluif.portOut[5]~51_combout ),
	.datac(\ShiftRight0~95_combout ),
	.datad(\ShiftRight0~92_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[5]~54_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~54 .lut_mask = 16'hE6A2;
defparam \aluif.portOut[5]~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N14
cycloneive_lcell_comb \aluif.portOut[5]~56 (
// Equation(s):
// \aluif.portOut[5]~56_combout  = (\aluif.portOut[5]~55_combout  & ((\prif.ALUOP_ex [2] & ((\aluif.portOut[5]~54_combout ))) # (!\prif.ALUOP_ex [2] & (\portOut~10_combout )))) # (!\aluif.portOut[5]~55_combout  & (!\prif.ALUOP_ex [2]))

	.dataa(\aluif.portOut[5]~55_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\portOut~10_combout ),
	.datad(\aluif.portOut[5]~54_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[5]~56_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~56 .lut_mask = 16'hB931;
defparam \aluif.portOut[5]~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N8
cycloneive_lcell_comb \Add0~8 (
// Equation(s):
// \Add0~8_combout  = ((\Mux27~1_combout  $ (\Mux91~2_combout  $ (!\Add0~7 )))) # (GND)
// \Add0~9  = CARRY((\Mux27~1_combout  & ((\Mux91~2_combout ) # (!\Add0~7 ))) # (!\Mux27~1_combout  & (\Mux91~2_combout  & !\Add0~7 )))

	.dataa(Mux27),
	.datab(Mux91),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~7 ),
	.combout(\Add0~8_combout ),
	.cout(\Add0~9 ));
// synopsys translate_off
defparam \Add0~8 .lut_mask = 16'h698E;
defparam \Add0~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N10
cycloneive_lcell_comb \Add0~10 (
// Equation(s):
// \Add0~10_combout  = (\Mux90~3_combout  & ((\Mux26~1_combout  & (\Add0~9  & VCC)) # (!\Mux26~1_combout  & (!\Add0~9 )))) # (!\Mux90~3_combout  & ((\Mux26~1_combout  & (!\Add0~9 )) # (!\Mux26~1_combout  & ((\Add0~9 ) # (GND)))))
// \Add0~11  = CARRY((\Mux90~3_combout  & (!\Mux26~1_combout  & !\Add0~9 )) # (!\Mux90~3_combout  & ((!\Add0~9 ) # (!\Mux26~1_combout ))))

	.dataa(Mux90),
	.datab(Mux26),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~9 ),
	.combout(\Add0~10_combout ),
	.cout(\Add0~11 ));
// synopsys translate_off
defparam \Add0~10 .lut_mask = 16'h9617;
defparam \Add0~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N8
cycloneive_lcell_comb \ShiftLeft0~18 (
// Equation(s):
// \ShiftLeft0~18_combout  = (\Mux95~1_combout  & ((\Mux29~1_combout ))) # (!\Mux95~1_combout  & (\Mux28~1_combout ))

	.dataa(Mux95),
	.datab(gnd),
	.datac(Mux28),
	.datad(Mux29),
	.cin(gnd),
	.combout(\ShiftLeft0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~18 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N12
cycloneive_lcell_comb \ShiftLeft0~23 (
// Equation(s):
// \ShiftLeft0~23_combout  = (\Mux95~1_combout  & ((\Mux27~1_combout ))) # (!\Mux95~1_combout  & (\Mux26~1_combout ))

	.dataa(Mux95),
	.datab(gnd),
	.datac(Mux26),
	.datad(Mux27),
	.cin(gnd),
	.combout(\ShiftLeft0~23_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~23 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N6
cycloneive_lcell_comb \ShiftLeft0~24 (
// Equation(s):
// \ShiftLeft0~24_combout  = (\Mux94~1_combout  & (\ShiftLeft0~18_combout )) # (!\Mux94~1_combout  & ((\ShiftLeft0~23_combout )))

	.dataa(Mux94),
	.datab(gnd),
	.datac(\ShiftLeft0~18_combout ),
	.datad(\ShiftLeft0~23_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~24_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~24 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y22_N24
cycloneive_lcell_comb \ShiftLeft0~22 (
// Equation(s):
// \ShiftLeft0~22_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux31~1_combout ))) # (!\Mux95~1_combout  & (\Mux30~1_combout ))))

	.dataa(Mux94),
	.datab(Mux95),
	.datac(Mux30),
	.datad(Mux31),
	.cin(gnd),
	.combout(\ShiftLeft0~22_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~22 .lut_mask = 16'h5410;
defparam \ShiftLeft0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y22_N10
cycloneive_lcell_comb \ShiftLeft0~25 (
// Equation(s):
// \ShiftLeft0~25_combout  = (!\Mux92~2_combout  & ((\Mux93~2_combout  & ((\ShiftLeft0~22_combout ))) # (!\Mux93~2_combout  & (\ShiftLeft0~24_combout ))))

	.dataa(Mux931),
	.datab(Mux92),
	.datac(\ShiftLeft0~24_combout ),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~25_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~25 .lut_mask = 16'h3210;
defparam \ShiftLeft0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N4
cycloneive_lcell_comb \aluif.portOut[5]~49 (
// Equation(s):
// \aluif.portOut[5]~49_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[15]~26_combout  & \ShiftLeft0~25_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~9_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(\portOut~9_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\ShiftLeft0~25_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[5]~49_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~49 .lut_mask = 16'hE323;
defparam \aluif.portOut[5]~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N24
cycloneive_lcell_comb \portOut~8 (
// Equation(s):
// \portOut~8_combout  = \Mux90~3_combout  $ (\Mux26~1_combout )

	.dataa(gnd),
	.datab(Mux90),
	.datac(gnd),
	.datad(Mux26),
	.cin(gnd),
	.combout(\portOut~8_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~8 .lut_mask = 16'h33CC;
defparam \portOut~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N30
cycloneive_lcell_comb \aluif.portOut[5]~50 (
// Equation(s):
// \aluif.portOut[5]~50_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[5]~49_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[5]~49_combout  & ((\portOut~8_combout ))) # (!\aluif.portOut[5]~49_combout  & (\Add0~10_combout ))))

	.dataa(prifALUOP_ex_1),
	.datab(\Add0~10_combout ),
	.datac(\aluif.portOut[5]~49_combout ),
	.datad(\portOut~8_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[5]~50_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~50 .lut_mask = 16'hF4A4;
defparam \aluif.portOut[5]~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N4
cycloneive_lcell_comb \portOut~11 (
// Equation(s):
// \portOut~11_combout  = \Mux27~1_combout  $ (\Mux91~2_combout )

	.dataa(Mux27),
	.datab(gnd),
	.datac(Mux91),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~11_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~11 .lut_mask = 16'h5A5A;
defparam \portOut~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N6
cycloneive_lcell_comb \portOut~12 (
// Equation(s):
// \portOut~12_combout  = (\Mux91~2_combout  & \Mux27~1_combout )

	.dataa(gnd),
	.datab(Mux91),
	.datac(gnd),
	.datad(Mux27),
	.cin(gnd),
	.combout(\portOut~12_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~12 .lut_mask = 16'hCC00;
defparam \portOut~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N28
cycloneive_lcell_comb \aluif.portOut[4]~59 (
// Equation(s):
// \aluif.portOut[4]~59_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & (\ShiftLeft0~29_combout )) # (!\prif.ALUOP_ex [2] & ((\portOut~12_combout ))))) # (!\aluif.portOut[15]~26_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\ShiftLeft0~29_combout ),
	.datab(\aluif.portOut[15]~26_combout ),
	.datac(prifALUOP_ex_2),
	.datad(\portOut~12_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[4]~59_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[4]~59 .lut_mask = 16'h8F83;
defparam \aluif.portOut[4]~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N14
cycloneive_lcell_comb \aluif.portOut[4]~60 (
// Equation(s):
// \aluif.portOut[4]~60_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[4]~59_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[4]~59_combout  & ((\portOut~11_combout ))) # (!\aluif.portOut[4]~59_combout  & (\Add0~8_combout ))))

	.dataa(\Add0~8_combout ),
	.datab(\portOut~11_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.portOut[4]~59_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[4]~60_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[4]~60 .lut_mask = 16'hFC0A;
defparam \aluif.portOut[4]~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N12
cycloneive_lcell_comb \portOut~13 (
// Equation(s):
// \portOut~13_combout  = (\Mux27~1_combout ) # (\Mux91~2_combout )

	.dataa(Mux27),
	.datab(gnd),
	.datac(Mux91),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~13_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~13 .lut_mask = 16'hFAFA;
defparam \portOut~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N30
cycloneive_lcell_comb \aluif.portOut[5]~52 (
// Equation(s):
// \aluif.portOut[5]~52_combout  = (\Mux91~2_combout ) # ((!\Mux92~2_combout  & \Mux93~2_combout ))

	.dataa(gnd),
	.datab(Mux92),
	.datac(Mux91),
	.datad(Mux931),
	.cin(gnd),
	.combout(\aluif.portOut[5]~52_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[5]~52 .lut_mask = 16'hF3F0;
defparam \aluif.portOut[5]~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N24
cycloneive_lcell_comb \aluif.portOut[4]~61 (
// Equation(s):
// \aluif.portOut[4]~61_combout  = (\aluif.portOut[5]~51_combout  & (((\aluif.portOut[5]~52_combout )))) # (!\aluif.portOut[5]~51_combout  & ((\aluif.portOut[5]~52_combout  & (\ShiftRight0~58_combout )) # (!\aluif.portOut[5]~52_combout  & 
// ((\ShiftRight0~51_combout )))))

	.dataa(\ShiftRight0~58_combout ),
	.datab(\aluif.portOut[5]~51_combout ),
	.datac(\aluif.portOut[5]~52_combout ),
	.datad(\ShiftRight0~51_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[4]~61_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[4]~61 .lut_mask = 16'hE3E0;
defparam \aluif.portOut[4]~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N6
cycloneive_lcell_comb \ShiftRight0~43 (
// Equation(s):
// \ShiftRight0~43_combout  = (\Mux95~1_combout  & (\Mux0~1_combout )) # (!\Mux95~1_combout  & ((\Mux1~1_combout )))

	.dataa(gnd),
	.datab(Mux95),
	.datac(Mux0),
	.datad(Mux1),
	.cin(gnd),
	.combout(\ShiftRight0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~43 .lut_mask = 16'hF3C0;
defparam \ShiftRight0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N24
cycloneive_lcell_comb \ShiftRight0~44 (
// Equation(s):
// \ShiftRight0~44_combout  = (\ShiftRight0~42_combout ) # ((\Mux94~1_combout  & \ShiftRight0~43_combout ))

	.dataa(\ShiftRight0~42_combout ),
	.datab(gnd),
	.datac(Mux94),
	.datad(\ShiftRight0~43_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~44 .lut_mask = 16'hFAAA;
defparam \ShiftRight0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N30
cycloneive_lcell_comb \ShiftRight0~98 (
// Equation(s):
// \ShiftRight0~98_combout  = (\Mux92~2_combout  & (((!\Mux93~2_combout  & \ShiftRight0~44_combout )))) # (!\Mux92~2_combout  & (\ShiftRight0~97_combout ))

	.dataa(\ShiftRight0~97_combout ),
	.datab(Mux931),
	.datac(Mux92),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~98 .lut_mask = 16'h3A0A;
defparam \ShiftRight0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N2
cycloneive_lcell_comb \aluif.portOut[4]~62 (
// Equation(s):
// \aluif.portOut[4]~62_combout  = (\aluif.portOut[4]~61_combout  & (((\ShiftRight0~98_combout ) # (!\aluif.portOut[5]~51_combout )))) # (!\aluif.portOut[4]~61_combout  & (\ShiftRight0~96_combout  & (\aluif.portOut[5]~51_combout )))

	.dataa(\ShiftRight0~96_combout ),
	.datab(\aluif.portOut[4]~61_combout ),
	.datac(\aluif.portOut[5]~51_combout ),
	.datad(\ShiftRight0~98_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[4]~62_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[4]~62 .lut_mask = 16'hEC2C;
defparam \aluif.portOut[4]~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N16
cycloneive_lcell_comb \aluif.portOut[4]~63 (
// Equation(s):
// \aluif.portOut[4]~63_combout  = (\aluif.portOut[5]~55_combout  & ((\prif.ALUOP_ex [2] & (\aluif.portOut[4]~62_combout )) # (!\prif.ALUOP_ex [2] & ((\portOut~13_combout ))))) # (!\aluif.portOut[5]~55_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\aluif.portOut[5]~55_combout ),
	.datab(\aluif.portOut[4]~62_combout ),
	.datac(prifALUOP_ex_2),
	.datad(\portOut~13_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[4]~63_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[4]~63 .lut_mask = 16'h8F85;
defparam \aluif.portOut[4]~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N30
cycloneive_lcell_comb \aluif.portOut[4]~64 (
// Equation(s):
// \aluif.portOut[4]~64_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[4]~63_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[4]~63_combout  & (!\portOut~13_combout )) # (!\aluif.portOut[4]~63_combout  & ((\Add1~8_combout )))))

	.dataa(\portOut~13_combout ),
	.datab(\Add1~8_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.portOut[4]~63_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[4]~64_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[4]~64 .lut_mask = 16'hF50C;
defparam \aluif.portOut[4]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N16
cycloneive_lcell_comb \ShiftRight0~75 (
// Equation(s):
// \ShiftRight0~75_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux13~1_combout )) # (!\Mux95~1_combout  & ((\Mux14~1_combout )))))

	.dataa(Mux94),
	.datab(Mux13),
	.datac(Mux95),
	.datad(Mux14),
	.cin(gnd),
	.combout(\ShiftRight0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~75 .lut_mask = 16'h8A80;
defparam \ShiftRight0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N22
cycloneive_lcell_comb \ShiftRight0~74 (
// Equation(s):
// \ShiftRight0~74_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux15~1_combout ))) # (!\Mux95~1_combout  & (\Mux16~1_combout ))))

	.dataa(Mux95),
	.datab(Mux16),
	.datac(Mux15),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftRight0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~74 .lut_mask = 16'h00E4;
defparam \ShiftRight0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N16
cycloneive_lcell_comb \ShiftRight0~68 (
// Equation(s):
// \ShiftRight0~68_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux9~1_combout ))) # (!\Mux95~1_combout  & (\Mux10~1_combout )))) # (!\Mux94~1_combout  & (\Mux95~1_combout ))

	.dataa(Mux94),
	.datab(Mux95),
	.datac(Mux10),
	.datad(Mux9),
	.cin(gnd),
	.combout(\ShiftRight0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~68 .lut_mask = 16'hEC64;
defparam \ShiftRight0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N10
cycloneive_lcell_comb \ShiftRight0~69 (
// Equation(s):
// \ShiftRight0~69_combout  = (\Mux94~1_combout  & (((\ShiftRight0~68_combout )))) # (!\Mux94~1_combout  & ((\ShiftRight0~68_combout  & ((\Mux11~1_combout ))) # (!\ShiftRight0~68_combout  & (\Mux12~1_combout ))))

	.dataa(Mux12),
	.datab(Mux11),
	.datac(Mux94),
	.datad(\ShiftRight0~68_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~69 .lut_mask = 16'hFC0A;
defparam \ShiftRight0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N24
cycloneive_lcell_comb \ShiftRight0~99 (
// Equation(s):
// \ShiftRight0~99_combout  = (\Mux93~2_combout  & (((\ShiftRight0~69_combout )))) # (!\Mux93~2_combout  & ((\ShiftRight0~75_combout ) # ((\ShiftRight0~74_combout ))))

	.dataa(Mux931),
	.datab(\ShiftRight0~75_combout ),
	.datac(\ShiftRight0~74_combout ),
	.datad(\ShiftRight0~69_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~99 .lut_mask = 16'hFE54;
defparam \ShiftRight0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N0
cycloneive_lcell_comb \aluif.portOut[7]~68 (
// Equation(s):
// \aluif.portOut[7]~68_combout  = (\aluif.portOut[5]~51_combout  & (((\ShiftRight0~99_combout ) # (\aluif.portOut[5]~52_combout )))) # (!\aluif.portOut[5]~51_combout  & (\ShiftRight0~72_combout  & ((!\aluif.portOut[5]~52_combout ))))

	.dataa(\ShiftRight0~72_combout ),
	.datab(\ShiftRight0~99_combout ),
	.datac(\aluif.portOut[5]~51_combout ),
	.datad(\aluif.portOut[5]~52_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[7]~68_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[7]~68 .lut_mask = 16'hF0CA;
defparam \aluif.portOut[7]~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N28
cycloneive_lcell_comb \ShiftRight0~16 (
// Equation(s):
// \ShiftRight0~16_combout  = (\Mux95~1_combout  & ((\Mux19~1_combout ) # ((\Mux19~0_combout )))) # (!\Mux95~1_combout  & (((\Mux20~1_combout ))))

	.dataa(Mux191),
	.datab(Mux19),
	.datac(Mux20),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~16_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~16 .lut_mask = 16'hEEF0;
defparam \ShiftRight0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N20
cycloneive_lcell_comb \ShiftRight0~73 (
// Equation(s):
// \ShiftRight0~73_combout  = (\Mux94~1_combout  & (\ShiftRight0~14_combout )) # (!\Mux94~1_combout  & ((\ShiftRight0~16_combout )))

	.dataa(Mux94),
	.datab(gnd),
	.datac(\ShiftRight0~14_combout ),
	.datad(\ShiftRight0~16_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~73 .lut_mask = 16'hF5A0;
defparam \ShiftRight0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N30
cycloneive_lcell_comb \ShiftRight0~64 (
// Equation(s):
// \ShiftRight0~64_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux3~1_combout ))) # (!\Mux95~1_combout  & (\Mux4~1_combout ))))

	.dataa(Mux95),
	.datab(Mux4),
	.datac(Mux3),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftRight0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~64 .lut_mask = 16'h00E4;
defparam \ShiftRight0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N2
cycloneive_lcell_comb \ShiftRight0~100 (
// Equation(s):
// \ShiftRight0~100_combout  = (\Mux93~2_combout  & ((\ShiftRight0~63_combout ) # ((\ShiftRight0~64_combout )))) # (!\Mux93~2_combout  & (((\ShiftRight0~67_combout ))))

	.dataa(Mux931),
	.datab(\ShiftRight0~63_combout ),
	.datac(\ShiftRight0~64_combout ),
	.datad(\ShiftRight0~67_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~100 .lut_mask = 16'hFDA8;
defparam \ShiftRight0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N28
cycloneive_lcell_comb \ShiftRight0~101 (
// Equation(s):
// \ShiftRight0~101_combout  = (\Mux92~2_combout  & (!\Mux93~2_combout  & (\ShiftRight0~62_combout ))) # (!\Mux92~2_combout  & (((\ShiftRight0~100_combout ))))

	.dataa(Mux931),
	.datab(\ShiftRight0~62_combout ),
	.datac(Mux92),
	.datad(\ShiftRight0~100_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~101 .lut_mask = 16'h4F40;
defparam \ShiftRight0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N22
cycloneive_lcell_comb \aluif.portOut[7]~69 (
// Equation(s):
// \aluif.portOut[7]~69_combout  = (\aluif.portOut[5]~52_combout  & ((\aluif.portOut[7]~68_combout  & ((\ShiftRight0~101_combout ))) # (!\aluif.portOut[7]~68_combout  & (\ShiftRight0~73_combout )))) # (!\aluif.portOut[5]~52_combout  & 
// (\aluif.portOut[7]~68_combout ))

	.dataa(\aluif.portOut[5]~52_combout ),
	.datab(\aluif.portOut[7]~68_combout ),
	.datac(\ShiftRight0~73_combout ),
	.datad(\ShiftRight0~101_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[7]~69_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[7]~69 .lut_mask = 16'hEC64;
defparam \aluif.portOut[7]~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N8
cycloneive_lcell_comb \aluif.portOut[7]~70 (
// Equation(s):
// \aluif.portOut[7]~70_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[7]~69_combout  & \aluif.portOut[5]~55_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~16_combout ) # ((!\aluif.portOut[5]~55_combout ))))

	.dataa(\portOut~16_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\aluif.portOut[7]~69_combout ),
	.datad(\aluif.portOut[5]~55_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[7]~70_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[7]~70 .lut_mask = 16'hE233;
defparam \aluif.portOut[7]~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N12
cycloneive_lcell_comb \Add1~12 (
// Equation(s):
// \Add1~12_combout  = ((\Mux25~1_combout  $ (\Mux89~4_combout  $ (\Add1~11 )))) # (GND)
// \Add1~13  = CARRY((\Mux25~1_combout  & ((!\Add1~11 ) # (!\Mux89~4_combout ))) # (!\Mux25~1_combout  & (!\Mux89~4_combout  & !\Add1~11 )))

	.dataa(Mux25),
	.datab(Mux891),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~11 ),
	.combout(\Add1~12_combout ),
	.cout(\Add1~13 ));
// synopsys translate_off
defparam \Add1~12 .lut_mask = 16'h962B;
defparam \Add1~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N14
cycloneive_lcell_comb \Add1~14 (
// Equation(s):
// \Add1~14_combout  = (\Mux24~1_combout  & ((\Mux88~3_combout  & (!\Add1~13 )) # (!\Mux88~3_combout  & (\Add1~13  & VCC)))) # (!\Mux24~1_combout  & ((\Mux88~3_combout  & ((\Add1~13 ) # (GND))) # (!\Mux88~3_combout  & (!\Add1~13 ))))
// \Add1~15  = CARRY((\Mux24~1_combout  & (\Mux88~3_combout  & !\Add1~13 )) # (!\Mux24~1_combout  & ((\Mux88~3_combout ) # (!\Add1~13 ))))

	.dataa(Mux24),
	.datab(Mux88),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~13 ),
	.combout(\Add1~14_combout ),
	.cout(\Add1~15 ));
// synopsys translate_off
defparam \Add1~14 .lut_mask = 16'h694D;
defparam \Add1~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N20
cycloneive_lcell_comb \portOut~16 (
// Equation(s):
// \portOut~16_combout  = (\Mux24~1_combout ) # (\Mux88~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux24),
	.datad(Mux88),
	.cin(gnd),
	.combout(\portOut~16_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~16 .lut_mask = 16'hFFF0;
defparam \portOut~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N26
cycloneive_lcell_comb \aluif.portOut[7]~71 (
// Equation(s):
// \aluif.portOut[7]~71_combout  = (\prif.ALUOP_ex [1] & (\aluif.portOut[7]~70_combout )) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[7]~70_combout  & ((!\portOut~16_combout ))) # (!\aluif.portOut[7]~70_combout  & (\Add1~14_combout ))))

	.dataa(prifALUOP_ex_1),
	.datab(\aluif.portOut[7]~70_combout ),
	.datac(\Add1~14_combout ),
	.datad(\portOut~16_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[7]~71_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[7]~71 .lut_mask = 16'h98DC;
defparam \aluif.portOut[7]~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N12
cycloneive_lcell_comb \Add0~12 (
// Equation(s):
// \Add0~12_combout  = ((\Mux25~1_combout  $ (\Mux89~4_combout  $ (!\Add0~11 )))) # (GND)
// \Add0~13  = CARRY((\Mux25~1_combout  & ((\Mux89~4_combout ) # (!\Add0~11 ))) # (!\Mux25~1_combout  & (\Mux89~4_combout  & !\Add0~11 )))

	.dataa(Mux25),
	.datab(Mux891),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~11 ),
	.combout(\Add0~12_combout ),
	.cout(\Add0~13 ));
// synopsys translate_off
defparam \Add0~12 .lut_mask = 16'h698E;
defparam \Add0~12 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N14
cycloneive_lcell_comb \Add0~14 (
// Equation(s):
// \Add0~14_combout  = (\Mux24~1_combout  & ((\Mux88~3_combout  & (\Add0~13  & VCC)) # (!\Mux88~3_combout  & (!\Add0~13 )))) # (!\Mux24~1_combout  & ((\Mux88~3_combout  & (!\Add0~13 )) # (!\Mux88~3_combout  & ((\Add0~13 ) # (GND)))))
// \Add0~15  = CARRY((\Mux24~1_combout  & (!\Mux88~3_combout  & !\Add0~13 )) # (!\Mux24~1_combout  & ((!\Add0~13 ) # (!\Mux88~3_combout ))))

	.dataa(Mux24),
	.datab(Mux88),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~13 ),
	.combout(\Add0~14_combout ),
	.cout(\Add0~15 ));
// synopsys translate_off
defparam \Add0~14 .lut_mask = 16'h9617;
defparam \Add0~14 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N28
cycloneive_lcell_comb \portOut~14 (
// Equation(s):
// \portOut~14_combout  = \Mux88~3_combout  $ (\Mux24~1_combout )

	.dataa(gnd),
	.datab(Mux88),
	.datac(gnd),
	.datad(Mux24),
	.cin(gnd),
	.combout(\portOut~14_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~14 .lut_mask = 16'h33CC;
defparam \portOut~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N18
cycloneive_lcell_comb \ShiftLeft0~31 (
// Equation(s):
// \ShiftLeft0~31_combout  = (\Mux95~1_combout  & ((\Mux25~1_combout ))) # (!\Mux95~1_combout  & (\Mux24~1_combout ))

	.dataa(Mux24),
	.datab(gnd),
	.datac(Mux25),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftLeft0~31_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~31 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N0
cycloneive_lcell_comb \ShiftLeft0~32 (
// Equation(s):
// \ShiftLeft0~32_combout  = (\Mux94~1_combout  & ((\ShiftLeft0~23_combout ))) # (!\Mux94~1_combout  & (\ShiftLeft0~31_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~31_combout ),
	.datac(Mux94),
	.datad(\ShiftLeft0~23_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~32_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~32 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N20
cycloneive_lcell_comb \ShiftLeft0~30 (
// Equation(s):
// \ShiftLeft0~30_combout  = (\Mux94~1_combout  & ((\ShiftLeft0~4_combout ))) # (!\Mux94~1_combout  & (\ShiftLeft0~18_combout ))

	.dataa(Mux94),
	.datab(gnd),
	.datac(\ShiftLeft0~18_combout ),
	.datad(\ShiftLeft0~4_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~30_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~30 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N24
cycloneive_lcell_comb \ShiftLeft0~33 (
// Equation(s):
// \ShiftLeft0~33_combout  = (!\Mux92~2_combout  & ((\Mux93~2_combout  & ((\ShiftLeft0~30_combout ))) # (!\Mux93~2_combout  & (\ShiftLeft0~32_combout ))))

	.dataa(Mux92),
	.datab(\ShiftLeft0~32_combout ),
	.datac(Mux931),
	.datad(\ShiftLeft0~30_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~33 .lut_mask = 16'h5404;
defparam \ShiftLeft0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N24
cycloneive_lcell_comb \aluif.portOut[7]~66 (
// Equation(s):
// \aluif.portOut[7]~66_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & ((\ShiftLeft0~33_combout ))) # (!\prif.ALUOP_ex [2] & (\portOut~15_combout )))) # (!\aluif.portOut[15]~26_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\portOut~15_combout ),
	.datab(\aluif.portOut[15]~26_combout ),
	.datac(\ShiftLeft0~33_combout ),
	.datad(prifALUOP_ex_2),
	.cin(gnd),
	.combout(\aluif.portOut[7]~66_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[7]~66 .lut_mask = 16'hC0BB;
defparam \aluif.portOut[7]~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N18
cycloneive_lcell_comb \aluif.portOut[7]~67 (
// Equation(s):
// \aluif.portOut[7]~67_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[7]~66_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[7]~66_combout  & ((\portOut~14_combout ))) # (!\aluif.portOut[7]~66_combout  & (\Add0~14_combout ))))

	.dataa(\Add0~14_combout ),
	.datab(\portOut~14_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.portOut[7]~66_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[7]~67_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[7]~67 .lut_mask = 16'hFC0A;
defparam \aluif.portOut[7]~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N18
cycloneive_lcell_comb \portOut~17 (
// Equation(s):
// \portOut~17_combout  = \Mux25~1_combout  $ (\Mux89~4_combout )

	.dataa(gnd),
	.datab(Mux25),
	.datac(Mux891),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~17_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~17 .lut_mask = 16'h3C3C;
defparam \portOut~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N20
cycloneive_lcell_comb \ShiftLeft0~34 (
// Equation(s):
// \ShiftLeft0~34_combout  = (\Mux95~1_combout  & (\Mux26~1_combout )) # (!\Mux95~1_combout  & ((\Mux25~1_combout )))

	.dataa(Mux26),
	.datab(gnd),
	.datac(Mux25),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftLeft0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~34 .lut_mask = 16'hAAF0;
defparam \ShiftLeft0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N30
cycloneive_lcell_comb \ShiftLeft0~35 (
// Equation(s):
// \ShiftLeft0~35_combout  = (\Mux94~1_combout  & (\ShiftLeft0~27_combout )) # (!\Mux94~1_combout  & ((\ShiftLeft0~34_combout )))

	.dataa(\ShiftLeft0~27_combout ),
	.datab(gnd),
	.datac(Mux94),
	.datad(\ShiftLeft0~34_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~35 .lut_mask = 16'hAFA0;
defparam \ShiftLeft0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N10
cycloneive_lcell_comb \ShiftLeft0~36 (
// Equation(s):
// \ShiftLeft0~36_combout  = (!\Mux92~2_combout  & ((\Mux93~2_combout  & (\ShiftLeft0~21_combout )) # (!\Mux93~2_combout  & ((\ShiftLeft0~35_combout )))))

	.dataa(Mux92),
	.datab(\ShiftLeft0~21_combout ),
	.datac(Mux931),
	.datad(\ShiftLeft0~35_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~36 .lut_mask = 16'h4540;
defparam \ShiftLeft0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N20
cycloneive_lcell_comb \portOut~18 (
// Equation(s):
// \portOut~18_combout  = (\Mux25~1_combout  & \Mux89~4_combout )

	.dataa(gnd),
	.datab(Mux25),
	.datac(Mux891),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~18_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~18 .lut_mask = 16'hC0C0;
defparam \portOut~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N2
cycloneive_lcell_comb \aluif.portOut[6]~73 (
// Equation(s):
// \aluif.portOut[6]~73_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & (\ShiftLeft0~36_combout )) # (!\prif.ALUOP_ex [2] & ((\portOut~18_combout ))))) # (!\aluif.portOut[15]~26_combout  & (!\prif.ALUOP_ex [2]))

	.dataa(\aluif.portOut[15]~26_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\ShiftLeft0~36_combout ),
	.datad(\portOut~18_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[6]~73_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[6]~73 .lut_mask = 16'hB391;
defparam \aluif.portOut[6]~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N8
cycloneive_lcell_comb \aluif.portOut[6]~74 (
// Equation(s):
// \aluif.portOut[6]~74_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[6]~73_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[6]~73_combout  & ((\portOut~17_combout ))) # (!\aluif.portOut[6]~73_combout  & (\Add0~12_combout ))))

	.dataa(\Add0~12_combout ),
	.datab(\portOut~17_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.portOut[6]~73_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[6]~74_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[6]~74 .lut_mask = 16'hFC0A;
defparam \aluif.portOut[6]~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N14
cycloneive_lcell_comb \portOut~19 (
// Equation(s):
// \portOut~19_combout  = (\Mux25~1_combout ) # (\Mux89~4_combout )

	.dataa(gnd),
	.datab(Mux25),
	.datac(Mux891),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~19_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~19 .lut_mask = 16'hFCFC;
defparam \portOut~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N16
cycloneive_lcell_comb \ShiftRight0~103 (
// Equation(s):
// \ShiftRight0~103_combout  = (\Mux93~2_combout  & (\ShiftRight0~79_combout )) # (!\Mux93~2_combout  & ((\ShiftRight0~82_combout )))

	.dataa(\ShiftRight0~79_combout ),
	.datab(gnd),
	.datac(Mux931),
	.datad(\ShiftRight0~82_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~103 .lut_mask = 16'hAFA0;
defparam \ShiftRight0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N30
cycloneive_lcell_comb \ShiftRight0~104 (
// Equation(s):
// \ShiftRight0~104_combout  = (\Mux92~2_combout  & (!\ShiftLeft0~5_combout  & ((\ShiftRight0~43_combout )))) # (!\Mux92~2_combout  & (((\ShiftRight0~103_combout ))))

	.dataa(\ShiftLeft0~5_combout ),
	.datab(Mux92),
	.datac(\ShiftRight0~103_combout ),
	.datad(\ShiftRight0~43_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~104 .lut_mask = 16'h7430;
defparam \ShiftRight0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N18
cycloneive_lcell_comb \ShiftRight0~83 (
// Equation(s):
// \ShiftRight0~83_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux10~1_combout ))) # (!\Mux95~1_combout  & (\Mux11~1_combout )))) # (!\Mux94~1_combout  & (((\Mux95~1_combout ))))

	.dataa(Mux94),
	.datab(Mux11),
	.datac(Mux10),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~83 .lut_mask = 16'hF588;
defparam \ShiftRight0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N4
cycloneive_lcell_comb \ShiftRight0~84 (
// Equation(s):
// \ShiftRight0~84_combout  = (\Mux94~1_combout  & (((\ShiftRight0~83_combout )))) # (!\Mux94~1_combout  & ((\ShiftRight0~83_combout  & (\Mux12~1_combout )) # (!\ShiftRight0~83_combout  & ((\Mux13~1_combout )))))

	.dataa(Mux94),
	.datab(Mux12),
	.datac(Mux13),
	.datad(\ShiftRight0~83_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~84 .lut_mask = 16'hEE50;
defparam \ShiftRight0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y21_N10
cycloneive_lcell_comb \ShiftRight0~102 (
// Equation(s):
// \ShiftRight0~102_combout  = (\Mux93~2_combout  & (((\ShiftRight0~84_combout )))) # (!\Mux93~2_combout  & ((\ShiftRight0~89_combout ) # ((\ShiftRight0~90_combout ))))

	.dataa(\ShiftRight0~89_combout ),
	.datab(\ShiftRight0~84_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~90_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~102 .lut_mask = 16'hCFCA;
defparam \ShiftRight0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N22
cycloneive_lcell_comb \aluif.portOut[6]~75 (
// Equation(s):
// \aluif.portOut[6]~75_combout  = (\aluif.portOut[5]~51_combout  & (((\aluif.portOut[5]~52_combout ) # (\ShiftRight0~102_combout )))) # (!\aluif.portOut[5]~51_combout  & (\ShiftRight0~87_combout  & (!\aluif.portOut[5]~52_combout )))

	.dataa(\ShiftRight0~87_combout ),
	.datab(\aluif.portOut[5]~51_combout ),
	.datac(\aluif.portOut[5]~52_combout ),
	.datad(\ShiftRight0~102_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[6]~75_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[6]~75 .lut_mask = 16'hCEC2;
defparam \aluif.portOut[6]~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N28
cycloneive_lcell_comb \aluif.portOut[6]~76 (
// Equation(s):
// \aluif.portOut[6]~76_combout  = (\aluif.portOut[5]~52_combout  & ((\aluif.portOut[6]~75_combout  & (\ShiftRight0~104_combout )) # (!\aluif.portOut[6]~75_combout  & ((\ShiftRight0~88_combout ))))) # (!\aluif.portOut[5]~52_combout  & 
// (((\aluif.portOut[6]~75_combout ))))

	.dataa(\aluif.portOut[5]~52_combout ),
	.datab(\ShiftRight0~104_combout ),
	.datac(\ShiftRight0~88_combout ),
	.datad(\aluif.portOut[6]~75_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[6]~76_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[6]~76 .lut_mask = 16'hDDA0;
defparam \aluif.portOut[6]~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N10
cycloneive_lcell_comb \aluif.portOut[6]~77 (
// Equation(s):
// \aluif.portOut[6]~77_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[5]~55_combout  & \aluif.portOut[6]~76_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~19_combout ) # ((!\aluif.portOut[5]~55_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\portOut~19_combout ),
	.datac(\aluif.portOut[5]~55_combout ),
	.datad(\aluif.portOut[6]~76_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[6]~77_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[6]~77 .lut_mask = 16'hE545;
defparam \aluif.portOut[6]~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y25_N0
cycloneive_lcell_comb \aluif.portOut[6]~78 (
// Equation(s):
// \aluif.portOut[6]~78_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[6]~77_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[6]~77_combout  & ((!\portOut~19_combout ))) # (!\aluif.portOut[6]~77_combout  & (\Add1~12_combout ))))

	.dataa(\Add1~12_combout ),
	.datab(\portOut~19_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.portOut[6]~77_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[6]~78_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[6]~78 .lut_mask = 16'hF30A;
defparam \aluif.portOut[6]~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N16
cycloneive_lcell_comb \Add1~16 (
// Equation(s):
// \Add1~16_combout  = ((\Mux87~3_combout  $ (\Mux23~1_combout  $ (\Add1~15 )))) # (GND)
// \Add1~17  = CARRY((\Mux87~3_combout  & (\Mux23~1_combout  & !\Add1~15 )) # (!\Mux87~3_combout  & ((\Mux23~1_combout ) # (!\Add1~15 ))))

	.dataa(Mux87),
	.datab(Mux23),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~15 ),
	.combout(\Add1~16_combout ),
	.cout(\Add1~17 ));
// synopsys translate_off
defparam \Add1~16 .lut_mask = 16'h964D;
defparam \Add1~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N18
cycloneive_lcell_comb \Add1~18 (
// Equation(s):
// \Add1~18_combout  = (\Mux22~1_combout  & ((\Mux86~3_combout  & (!\Add1~17 )) # (!\Mux86~3_combout  & (\Add1~17  & VCC)))) # (!\Mux22~1_combout  & ((\Mux86~3_combout  & ((\Add1~17 ) # (GND))) # (!\Mux86~3_combout  & (!\Add1~17 ))))
// \Add1~19  = CARRY((\Mux22~1_combout  & (\Mux86~3_combout  & !\Add1~17 )) # (!\Mux22~1_combout  & ((\Mux86~3_combout ) # (!\Add1~17 ))))

	.dataa(Mux22),
	.datab(Mux86),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~17 ),
	.combout(\Add1~18_combout ),
	.cout(\Add1~19 ));
// synopsys translate_off
defparam \Add1~18 .lut_mask = 16'h694D;
defparam \Add1~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N20
cycloneive_lcell_comb \aluif.portOut[15]~80 (
// Equation(s):
// \aluif.portOut[15]~80_combout  = (!\prif.ALUOP_ex [1] & !\prif.ALUOP_ex [0])

	.dataa(gnd),
	.datab(gnd),
	.datac(prifALUOP_ex_1),
	.datad(prifALUOP_ex_0),
	.cin(gnd),
	.combout(\aluif.portOut[15]~80_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~80 .lut_mask = 16'h000F;
defparam \aluif.portOut[15]~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N28
cycloneive_lcell_comb \ShiftRight0~18 (
// Equation(s):
// \ShiftRight0~18_combout  = (\Mux94~1_combout  & (\ShiftRight0~16_combout )) # (!\Mux94~1_combout  & ((\ShiftRight0~17_combout )))

	.dataa(\ShiftRight0~16_combout ),
	.datab(\ShiftRight0~17_combout ),
	.datac(Mux94),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~18_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~18 .lut_mask = 16'hACAC;
defparam \ShiftRight0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y21_N10
cycloneive_lcell_comb \ShiftRight0~19 (
// Equation(s):
// \ShiftRight0~19_combout  = (\Mux93~2_combout  & ((\ShiftRight0~15_combout ))) # (!\Mux93~2_combout  & (\ShiftRight0~18_combout ))

	.dataa(gnd),
	.datab(\ShiftRight0~18_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~15_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~19 .lut_mask = 16'hFC0C;
defparam \ShiftRight0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N0
cycloneive_lcell_comb \aluif.portOut[15]~81 (
// Equation(s):
// \aluif.portOut[15]~81_combout  = ((\ShiftLeft0~15_combout ) # (\Mux91~2_combout )) # (!\prif.ALUOP_ex [2])

	.dataa(prifALUOP_ex_2),
	.datab(gnd),
	.datac(\ShiftLeft0~15_combout ),
	.datad(Mux91),
	.cin(gnd),
	.combout(\aluif.portOut[15]~81_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~81 .lut_mask = 16'hFFF5;
defparam \aluif.portOut[15]~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N8
cycloneive_lcell_comb \aluif.portOut[9]~85 (
// Equation(s):
// \aluif.portOut[9]~85_combout  = (\aluif.portOut[9]~84_combout  & (((\ShiftRight0~25_combout ) # (\aluif.portOut[15]~81_combout )))) # (!\aluif.portOut[9]~84_combout  & (\ShiftRight0~19_combout  & ((!\aluif.portOut[15]~81_combout ))))

	.dataa(\aluif.portOut[9]~84_combout ),
	.datab(\ShiftRight0~19_combout ),
	.datac(\ShiftRight0~25_combout ),
	.datad(\aluif.portOut[15]~81_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[9]~85_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[9]~85 .lut_mask = 16'hAAE4;
defparam \aluif.portOut[9]~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N22
cycloneive_lcell_comb \aluif.portOut[15]~86 (
// Equation(s):
// \aluif.portOut[15]~86_combout  = (!\prif.ALUOP_ex [0] & ((\prif.ALUOP_ex [1]) # (!\prif.ALUOP_ex [2])))

	.dataa(prifALUOP_ex_2),
	.datab(gnd),
	.datac(prifALUOP_ex_1),
	.datad(prifALUOP_ex_0),
	.cin(gnd),
	.combout(\aluif.portOut[15]~86_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~86 .lut_mask = 16'h00F5;
defparam \aluif.portOut[15]~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y21_N4
cycloneive_lcell_comb \portOut~21 (
// Equation(s):
// \portOut~21_combout  = \Mux86~3_combout  $ (\Mux22~1_combout )

	.dataa(gnd),
	.datab(Mux86),
	.datac(gnd),
	.datad(Mux22),
	.cin(gnd),
	.combout(\portOut~21_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~21 .lut_mask = 16'h33CC;
defparam \portOut~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N16
cycloneive_lcell_comb \Add0~16 (
// Equation(s):
// \Add0~16_combout  = ((\Mux23~1_combout  $ (\Mux87~3_combout  $ (!\Add0~15 )))) # (GND)
// \Add0~17  = CARRY((\Mux23~1_combout  & ((\Mux87~3_combout ) # (!\Add0~15 ))) # (!\Mux23~1_combout  & (\Mux87~3_combout  & !\Add0~15 )))

	.dataa(Mux23),
	.datab(Mux87),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~15 ),
	.combout(\Add0~16_combout ),
	.cout(\Add0~17 ));
// synopsys translate_off
defparam \Add0~16 .lut_mask = 16'h698E;
defparam \Add0~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N18
cycloneive_lcell_comb \Add0~18 (
// Equation(s):
// \Add0~18_combout  = (\Mux86~3_combout  & ((\Mux22~1_combout  & (\Add0~17  & VCC)) # (!\Mux22~1_combout  & (!\Add0~17 )))) # (!\Mux86~3_combout  & ((\Mux22~1_combout  & (!\Add0~17 )) # (!\Mux22~1_combout  & ((\Add0~17 ) # (GND)))))
// \Add0~19  = CARRY((\Mux86~3_combout  & (!\Mux22~1_combout  & !\Add0~17 )) # (!\Mux86~3_combout  & ((!\Add0~17 ) # (!\Mux22~1_combout ))))

	.dataa(Mux86),
	.datab(Mux22),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~17 ),
	.combout(\Add0~18_combout ),
	.cout(\Add0~19 ));
// synopsys translate_off
defparam \Add0~18 .lut_mask = 16'h9617;
defparam \Add0~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X57_Y21_N2
cycloneive_lcell_comb \portOut~22 (
// Equation(s):
// \portOut~22_combout  = (\Mux86~3_combout  & \Mux22~1_combout )

	.dataa(gnd),
	.datab(Mux86),
	.datac(gnd),
	.datad(Mux22),
	.cin(gnd),
	.combout(\portOut~22_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~22 .lut_mask = 16'hCC00;
defparam \portOut~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N0
cycloneive_lcell_comb \ShiftLeft0~37 (
// Equation(s):
// \ShiftLeft0~37_combout  = (\Mux95~1_combout  & (\Mux23~1_combout )) # (!\Mux95~1_combout  & ((\Mux22~1_combout )))

	.dataa(gnd),
	.datab(Mux23),
	.datac(Mux95),
	.datad(Mux22),
	.cin(gnd),
	.combout(\ShiftLeft0~37_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~37 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N14
cycloneive_lcell_comb \ShiftLeft0~38 (
// Equation(s):
// \ShiftLeft0~38_combout  = (\Mux94~1_combout  & ((\ShiftLeft0~31_combout ))) # (!\Mux94~1_combout  & (\ShiftLeft0~37_combout ))

	.dataa(Mux94),
	.datab(gnd),
	.datac(\ShiftLeft0~37_combout ),
	.datad(\ShiftLeft0~31_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~38 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N4
cycloneive_lcell_comb \ShiftLeft0~39 (
// Equation(s):
// \ShiftLeft0~39_combout  = (\Mux93~2_combout  & ((\ShiftLeft0~24_combout ))) # (!\Mux93~2_combout  & (\ShiftLeft0~38_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~38_combout ),
	.datac(Mux931),
	.datad(\ShiftLeft0~24_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~39 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N2
cycloneive_lcell_comb \ShiftLeft0~40 (
// Equation(s):
// \ShiftLeft0~40_combout  = (\Mux92~2_combout  & (\ShiftLeft0~4_combout  & ((!\ShiftLeft0~5_combout )))) # (!\Mux92~2_combout  & (((\ShiftLeft0~39_combout ))))

	.dataa(\ShiftLeft0~4_combout ),
	.datab(Mux92),
	.datac(\ShiftLeft0~39_combout ),
	.datad(\ShiftLeft0~5_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~40 .lut_mask = 16'h30B8;
defparam \ShiftLeft0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y21_N12
cycloneive_lcell_comb \aluif.portOut[9]~87 (
// Equation(s):
// \aluif.portOut[9]~87_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[15]~26_combout  & \ShiftLeft0~40_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~22_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\portOut~22_combout ),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\ShiftLeft0~40_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[9]~87_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[9]~87 .lut_mask = 16'hE545;
defparam \aluif.portOut[9]~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y21_N22
cycloneive_lcell_comb \aluif.portOut[9]~88 (
// Equation(s):
// \aluif.portOut[9]~88_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[9]~87_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[9]~87_combout  & (\portOut~21_combout )) # (!\aluif.portOut[9]~87_combout  & ((\Add0~18_combout )))))

	.dataa(prifALUOP_ex_1),
	.datab(\portOut~21_combout ),
	.datac(\Add0~18_combout ),
	.datad(\aluif.portOut[9]~87_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[9]~88_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[9]~88 .lut_mask = 16'hEE50;
defparam \aluif.portOut[9]~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N30
cycloneive_lcell_comb \aluif.portOut[9]~89 (
// Equation(s):
// \aluif.portOut[9]~89_combout  = (\aluif.portOut[15]~80_combout  & (((\aluif.portOut[15]~86_combout )))) # (!\aluif.portOut[15]~80_combout  & ((\aluif.portOut[15]~86_combout  & (\aluif.portOut[9]~85_combout )) # (!\aluif.portOut[15]~86_combout  & 
// ((\aluif.portOut[9]~88_combout )))))

	.dataa(\aluif.portOut[9]~85_combout ),
	.datab(\aluif.portOut[15]~80_combout ),
	.datac(\aluif.portOut[15]~86_combout ),
	.datad(\aluif.portOut[9]~88_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[9]~89_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[9]~89 .lut_mask = 16'hE3E0;
defparam \aluif.portOut[9]~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N16
cycloneive_lcell_comb \portOut~20 (
// Equation(s):
// \portOut~20_combout  = (\Mux22~1_combout ) # (\Mux86~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux22),
	.datad(Mux86),
	.cin(gnd),
	.combout(\portOut~20_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~20 .lut_mask = 16'hFFF0;
defparam \portOut~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N22
cycloneive_lcell_comb \portOut~23 (
// Equation(s):
// \portOut~23_combout  = (\Mux23~1_combout ) # (\Mux87~3_combout )

	.dataa(Mux23),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux87),
	.cin(gnd),
	.combout(\portOut~23_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~23 .lut_mask = 16'hFFAA;
defparam \portOut~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N20
cycloneive_lcell_comb \portOut~24 (
// Equation(s):
// \portOut~24_combout  = \Mux23~1_combout  $ (\Mux87~3_combout )

	.dataa(Mux23),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux87),
	.cin(gnd),
	.combout(\portOut~24_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~24 .lut_mask = 16'h55AA;
defparam \portOut~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N2
cycloneive_lcell_comb \ShiftLeft0~110 (
// Equation(s):
// \ShiftLeft0~110_combout  = (\Mux31~1_combout  & (!\Mux94~1_combout  & !\Mux95~1_combout ))

	.dataa(Mux31),
	.datab(Mux94),
	.datac(gnd),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftLeft0~110_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~110 .lut_mask = 16'h0022;
defparam \ShiftLeft0~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N28
cycloneive_lcell_comb \ShiftLeft0~26 (
// Equation(s):
// \ShiftLeft0~26_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux30~1_combout ))) # (!\Mux95~1_combout  & (\Mux29~1_combout ))))

	.dataa(Mux29),
	.datab(Mux94),
	.datac(Mux30),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftLeft0~26_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~26 .lut_mask = 16'hC088;
defparam \ShiftLeft0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N8
cycloneive_lcell_comb \ShiftLeft0~28 (
// Equation(s):
// \ShiftLeft0~28_combout  = (\ShiftLeft0~26_combout ) # ((\ShiftLeft0~27_combout  & !\Mux94~1_combout ))

	.dataa(\ShiftLeft0~27_combout ),
	.datab(gnd),
	.datac(Mux94),
	.datad(\ShiftLeft0~26_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~28_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~28 .lut_mask = 16'hFF0A;
defparam \ShiftLeft0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N0
cycloneive_lcell_comb \ShiftLeft0~41 (
// Equation(s):
// \ShiftLeft0~41_combout  = (\Mux95~1_combout  & ((\Mux24~1_combout ))) # (!\Mux95~1_combout  & (\Mux23~1_combout ))

	.dataa(gnd),
	.datab(Mux95),
	.datac(Mux23),
	.datad(Mux24),
	.cin(gnd),
	.combout(\ShiftLeft0~41_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~41 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N18
cycloneive_lcell_comb \ShiftLeft0~42 (
// Equation(s):
// \ShiftLeft0~42_combout  = (\Mux94~1_combout  & ((\ShiftLeft0~34_combout ))) # (!\Mux94~1_combout  & (\ShiftLeft0~41_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~41_combout ),
	.datac(Mux94),
	.datad(\ShiftLeft0~34_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~42 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N12
cycloneive_lcell_comb \ShiftLeft0~43 (
// Equation(s):
// \ShiftLeft0~43_combout  = (\Mux93~2_combout  & (\ShiftLeft0~28_combout )) # (!\Mux93~2_combout  & ((\ShiftLeft0~42_combout )))

	.dataa(Mux931),
	.datab(gnd),
	.datac(\ShiftLeft0~28_combout ),
	.datad(\ShiftLeft0~42_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~43_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~43 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N26
cycloneive_lcell_comb \ShiftLeft0~44 (
// Equation(s):
// \ShiftLeft0~44_combout  = (\Mux92~2_combout  & (!\Mux93~2_combout  & (\ShiftLeft0~110_combout ))) # (!\Mux92~2_combout  & (((\ShiftLeft0~43_combout ))))

	.dataa(Mux931),
	.datab(\ShiftLeft0~110_combout ),
	.datac(Mux92),
	.datad(\ShiftLeft0~43_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~44_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~44 .lut_mask = 16'h4F40;
defparam \ShiftLeft0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N12
cycloneive_lcell_comb \aluif.portOut[8]~93 (
// Equation(s):
// \aluif.portOut[8]~93_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & ((\ShiftLeft0~44_combout ))) # (!\prif.ALUOP_ex [2] & (\portOut~25_combout )))) # (!\aluif.portOut[15]~26_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\portOut~25_combout ),
	.datab(\ShiftLeft0~44_combout ),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(prifALUOP_ex_2),
	.cin(gnd),
	.combout(\aluif.portOut[8]~93_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[8]~93 .lut_mask = 16'hC0AF;
defparam \aluif.portOut[8]~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N6
cycloneive_lcell_comb \aluif.portOut[8]~94 (
// Equation(s):
// \aluif.portOut[8]~94_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[8]~93_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[8]~93_combout  & (\portOut~24_combout )) # (!\aluif.portOut[8]~93_combout  & ((\Add0~16_combout )))))

	.dataa(prifALUOP_ex_1),
	.datab(\portOut~24_combout ),
	.datac(\Add0~16_combout ),
	.datad(\aluif.portOut[8]~93_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[8]~94_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[8]~94 .lut_mask = 16'hEE50;
defparam \aluif.portOut[8]~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N0
cycloneive_lcell_comb \aluif.portOut[8]~95 (
// Equation(s):
// \aluif.portOut[8]~95_combout  = (\aluif.portOut[15]~86_combout  & (\aluif.portOut[15]~80_combout )) # (!\aluif.portOut[15]~86_combout  & ((\aluif.portOut[15]~80_combout  & (\Add1~16_combout )) # (!\aluif.portOut[15]~80_combout  & 
// ((\aluif.portOut[8]~94_combout )))))

	.dataa(\aluif.portOut[15]~86_combout ),
	.datab(\aluif.portOut[15]~80_combout ),
	.datac(\Add1~16_combout ),
	.datad(\aluif.portOut[8]~94_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[8]~95_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[8]~95 .lut_mask = 16'hD9C8;
defparam \aluif.portOut[8]~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N0
cycloneive_lcell_comb \ShiftRight0~36 (
// Equation(s):
// \ShiftRight0~36_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux10~1_combout ))) # (!\Mux95~1_combout  & (\Mux11~1_combout ))))

	.dataa(Mux95),
	.datab(Mux11),
	.datac(Mux10),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftRight0~36_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~36 .lut_mask = 16'h00E4;
defparam \ShiftRight0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N28
cycloneive_lcell_comb \ShiftRight0~34 (
// Equation(s):
// \ShiftRight0~34_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux12~1_combout )) # (!\Mux95~1_combout  & ((\Mux13~1_combout )))))

	.dataa(Mux95),
	.datab(Mux94),
	.datac(Mux12),
	.datad(Mux13),
	.cin(gnd),
	.combout(\ShiftRight0~34_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~34 .lut_mask = 16'hC480;
defparam \ShiftRight0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N10
cycloneive_lcell_comb \ShiftRight0~33 (
// Equation(s):
// \ShiftRight0~33_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux14~1_combout ))) # (!\Mux95~1_combout  & (\Mux15~1_combout ))))

	.dataa(Mux15),
	.datab(Mux94),
	.datac(Mux14),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~33_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~33 .lut_mask = 16'h3022;
defparam \ShiftRight0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N18
cycloneive_lcell_comb \ShiftRight0~35 (
// Equation(s):
// \ShiftRight0~35_combout  = (\ShiftRight0~34_combout ) # (\ShiftRight0~33_combout )

	.dataa(gnd),
	.datab(\ShiftRight0~34_combout ),
	.datac(gnd),
	.datad(\ShiftRight0~33_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~35_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~35 .lut_mask = 16'hFFCC;
defparam \ShiftRight0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N20
cycloneive_lcell_comb \ShiftRight0~38 (
// Equation(s):
// \ShiftRight0~38_combout  = (\Mux93~2_combout  & ((\ShiftRight0~37_combout ) # ((\ShiftRight0~36_combout )))) # (!\Mux93~2_combout  & (((\ShiftRight0~35_combout ))))

	.dataa(\ShiftRight0~37_combout ),
	.datab(\ShiftRight0~36_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~35_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~38_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~38 .lut_mask = 16'hEFE0;
defparam \ShiftRight0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N4
cycloneive_lcell_comb \ShiftRight0~106 (
// Equation(s):
// \ShiftRight0~106_combout  = (!\Mux92~2_combout  & ((\Mux93~2_combout  & ((\ShiftRight0~44_combout ))) # (!\Mux93~2_combout  & (\ShiftRight0~40_combout ))))

	.dataa(\ShiftRight0~40_combout ),
	.datab(Mux931),
	.datac(Mux92),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~106_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~106 .lut_mask = 16'h0E02;
defparam \ShiftRight0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N18
cycloneive_lcell_comb \aluif.portOut[15]~82 (
// Equation(s):
// \aluif.portOut[15]~82_combout  = ((\Mux91~2_combout  & !\ShiftLeft0~15_combout )) # (!\prif.ALUOP_ex [2])

	.dataa(gnd),
	.datab(Mux91),
	.datac(prifALUOP_ex_2),
	.datad(\ShiftLeft0~15_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[15]~82_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~82 .lut_mask = 16'h0FCF;
defparam \aluif.portOut[15]~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N20
cycloneive_lcell_comb \aluif.portOut[15]~83 (
// Equation(s):
// \aluif.portOut[15]~83_combout  = ((\Mux92~2_combout  & (!\Mux91~2_combout  & !\ShiftLeft0~15_combout ))) # (!\prif.ALUOP_ex [2])

	.dataa(Mux92),
	.datab(Mux91),
	.datac(prifALUOP_ex_2),
	.datad(\ShiftLeft0~15_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[15]~83_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~83 .lut_mask = 16'h0F2F;
defparam \aluif.portOut[15]~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N28
cycloneive_lcell_comb \aluif.portOut[8]~91 (
// Equation(s):
// \aluif.portOut[8]~91_combout  = (\aluif.portOut[15]~82_combout  & ((\aluif.portOut[15]~83_combout  & (\portOut~23_combout )) # (!\aluif.portOut[15]~83_combout  & ((\ShiftRight0~106_combout ))))) # (!\aluif.portOut[15]~82_combout  & 
// (((\aluif.portOut[15]~83_combout ))))

	.dataa(\portOut~23_combout ),
	.datab(\ShiftRight0~106_combout ),
	.datac(\aluif.portOut[15]~82_combout ),
	.datad(\aluif.portOut[15]~83_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[8]~91_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[8]~91 .lut_mask = 16'hAFC0;
defparam \aluif.portOut[8]~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N26
cycloneive_lcell_comb \aluif.portOut[8]~92 (
// Equation(s):
// \aluif.portOut[8]~92_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[8]~91_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[8]~91_combout  & ((\ShiftRight0~38_combout ))) # (!\aluif.portOut[8]~91_combout  & 
// (\ShiftRight0~59_combout ))))

	.dataa(\ShiftRight0~59_combout ),
	.datab(\aluif.portOut[15]~81_combout ),
	.datac(\ShiftRight0~38_combout ),
	.datad(\aluif.portOut[8]~91_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[8]~92_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[8]~92 .lut_mask = 16'hFC22;
defparam \aluif.portOut[8]~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N30
cycloneive_lcell_comb \portOut~26 (
// Equation(s):
// \portOut~26_combout  = (\Mux20~1_combout ) # (\Mux84~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux20),
	.datad(Mux84),
	.cin(gnd),
	.combout(\portOut~26_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~26 .lut_mask = 16'hFFF0;
defparam \portOut~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N26
cycloneive_lcell_comb \ShiftRight0~76 (
// Equation(s):
// \ShiftRight0~76_combout  = (\Mux93~2_combout  & (((\ShiftRight0~74_combout ) # (\ShiftRight0~75_combout )))) # (!\Mux93~2_combout  & (\ShiftRight0~73_combout ))

	.dataa(Mux931),
	.datab(\ShiftRight0~73_combout ),
	.datac(\ShiftRight0~74_combout ),
	.datad(\ShiftRight0~75_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~76 .lut_mask = 16'hEEE4;
defparam \ShiftRight0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N18
cycloneive_lcell_comb \ShiftRight0~107 (
// Equation(s):
// \ShiftRight0~107_combout  = (!\Mux92~2_combout  & \ShiftRight0~65_combout )

	.dataa(gnd),
	.datab(Mux92),
	.datac(\ShiftRight0~65_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\ShiftRight0~107_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~107 .lut_mask = 16'h3030;
defparam \ShiftRight0~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N12
cycloneive_lcell_comb \aluif.portOut[11]~97 (
// Equation(s):
// \aluif.portOut[11]~97_combout  = (\aluif.portOut[15]~83_combout  & (((\portOut~26_combout ) # (!\aluif.portOut[15]~82_combout )))) # (!\aluif.portOut[15]~83_combout  & (\ShiftRight0~107_combout  & ((\aluif.portOut[15]~82_combout ))))

	.dataa(\aluif.portOut[15]~83_combout ),
	.datab(\ShiftRight0~107_combout ),
	.datac(\portOut~26_combout ),
	.datad(\aluif.portOut[15]~82_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[11]~97_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[11]~97 .lut_mask = 16'hE4AA;
defparam \aluif.portOut[11]~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N14
cycloneive_lcell_comb \aluif.portOut[11]~98 (
// Equation(s):
// \aluif.portOut[11]~98_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[11]~97_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[11]~97_combout  & (\ShiftRight0~70_combout )) # (!\aluif.portOut[11]~97_combout  & 
// ((\ShiftRight0~76_combout )))))

	.dataa(\ShiftRight0~70_combout ),
	.datab(\aluif.portOut[15]~81_combout ),
	.datac(\ShiftRight0~76_combout ),
	.datad(\aluif.portOut[11]~97_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[11]~98_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[11]~98 .lut_mask = 16'hEE30;
defparam \aluif.portOut[11]~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N0
cycloneive_lcell_comb \portOut~27 (
// Equation(s):
// \portOut~27_combout  = \Mux20~1_combout  $ (\Mux84~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux20),
	.datad(Mux84),
	.cin(gnd),
	.combout(\portOut~27_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~27 .lut_mask = 16'h0FF0;
defparam \portOut~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N8
cycloneive_lcell_comb \ShiftLeft0~46 (
// Equation(s):
// \ShiftLeft0~46_combout  = (\Mux94~1_combout  & ((\ShiftLeft0~37_combout ))) # (!\Mux94~1_combout  & (\ShiftLeft0~45_combout ))

	.dataa(\ShiftLeft0~45_combout ),
	.datab(gnd),
	.datac(Mux94),
	.datad(\ShiftLeft0~37_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~46_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~46 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N28
cycloneive_lcell_comb \ShiftLeft0~47 (
// Equation(s):
// \ShiftLeft0~47_combout  = (\Mux93~2_combout  & ((\ShiftLeft0~32_combout ))) # (!\Mux93~2_combout  & (\ShiftLeft0~46_combout ))

	.dataa(Mux931),
	.datab(gnd),
	.datac(\ShiftLeft0~46_combout ),
	.datad(\ShiftLeft0~32_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~47_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~47 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N22
cycloneive_lcell_comb \ShiftLeft0~48 (
// Equation(s):
// \ShiftLeft0~48_combout  = (\Mux92~2_combout  & (\ShiftLeft0~30_combout  & (!\Mux93~2_combout ))) # (!\Mux92~2_combout  & (((\ShiftLeft0~47_combout ))))

	.dataa(Mux92),
	.datab(\ShiftLeft0~30_combout ),
	.datac(Mux931),
	.datad(\ShiftLeft0~47_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~48_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~48 .lut_mask = 16'h5D08;
defparam \ShiftLeft0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N28
cycloneive_lcell_comb \aluif.portOut[11]~99 (
// Equation(s):
// \aluif.portOut[11]~99_combout  = (\prif.ALUOP_ex [2] & (((\ShiftLeft0~48_combout  & \aluif.portOut[15]~26_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~28_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(\portOut~28_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\ShiftLeft0~48_combout ),
	.datad(\aluif.portOut[15]~26_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[11]~99_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[11]~99 .lut_mask = 16'hE233;
defparam \aluif.portOut[11]~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N2
cycloneive_lcell_comb \aluif.portOut[11]~100 (
// Equation(s):
// \aluif.portOut[11]~100_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[11]~99_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[11]~99_combout  & ((\portOut~27_combout ))) # (!\aluif.portOut[11]~99_combout  & (\Add0~22_combout ))))

	.dataa(\Add0~22_combout ),
	.datab(\portOut~27_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.portOut[11]~99_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[11]~100_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[11]~100 .lut_mask = 16'hFC0A;
defparam \aluif.portOut[11]~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y24_N0
cycloneive_lcell_comb \aluif.portOut[11]~101 (
// Equation(s):
// \aluif.portOut[11]~101_combout  = (\aluif.portOut[15]~86_combout  & ((\aluif.portOut[15]~80_combout ) # ((\aluif.portOut[11]~98_combout )))) # (!\aluif.portOut[15]~86_combout  & (!\aluif.portOut[15]~80_combout  & ((\aluif.portOut[11]~100_combout ))))

	.dataa(\aluif.portOut[15]~86_combout ),
	.datab(\aluif.portOut[15]~80_combout ),
	.datac(\aluif.portOut[11]~98_combout ),
	.datad(\aluif.portOut[11]~100_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[11]~101_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[11]~101 .lut_mask = 16'hB9A8;
defparam \aluif.portOut[11]~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N20
cycloneive_lcell_comb \Add1~20 (
// Equation(s):
// \Add1~20_combout  = ((\Mux21~1_combout  $ (\Mux85~3_combout  $ (\Add1~19 )))) # (GND)
// \Add1~21  = CARRY((\Mux21~1_combout  & ((!\Add1~19 ) # (!\Mux85~3_combout ))) # (!\Mux21~1_combout  & (!\Mux85~3_combout  & !\Add1~19 )))

	.dataa(Mux21),
	.datab(Mux85),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~19 ),
	.combout(\Add1~20_combout ),
	.cout(\Add1~21 ));
// synopsys translate_off
defparam \Add1~20 .lut_mask = 16'h962B;
defparam \Add1~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N22
cycloneive_lcell_comb \Add1~22 (
// Equation(s):
// \Add1~22_combout  = (\Mux84~3_combout  & ((\Mux20~1_combout  & (!\Add1~21 )) # (!\Mux20~1_combout  & ((\Add1~21 ) # (GND))))) # (!\Mux84~3_combout  & ((\Mux20~1_combout  & (\Add1~21  & VCC)) # (!\Mux20~1_combout  & (!\Add1~21 ))))
// \Add1~23  = CARRY((\Mux84~3_combout  & ((!\Add1~21 ) # (!\Mux20~1_combout ))) # (!\Mux84~3_combout  & (!\Mux20~1_combout  & !\Add1~21 )))

	.dataa(Mux84),
	.datab(Mux20),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~21 ),
	.combout(\Add1~22_combout ),
	.cout(\Add1~23 ));
// synopsys translate_off
defparam \Add1~22 .lut_mask = 16'h692B;
defparam \Add1~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N22
cycloneive_lcell_comb \portOut~29 (
// Equation(s):
// \portOut~29_combout  = (\Mux21~1_combout ) # (\Mux85~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux21),
	.datad(Mux85),
	.cin(gnd),
	.combout(\portOut~29_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~29 .lut_mask = 16'hFFF0;
defparam \portOut~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N8
cycloneive_lcell_comb \portOut~30 (
// Equation(s):
// \portOut~30_combout  = \Mux21~1_combout  $ (\Mux85~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux21),
	.datad(Mux85),
	.cin(gnd),
	.combout(\portOut~30_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~30 .lut_mask = 16'h0FF0;
defparam \portOut~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N20
cycloneive_lcell_comb \Add0~20 (
// Equation(s):
// \Add0~20_combout  = ((\Mux21~1_combout  $ (\Mux85~3_combout  $ (!\Add0~19 )))) # (GND)
// \Add0~21  = CARRY((\Mux21~1_combout  & ((\Mux85~3_combout ) # (!\Add0~19 ))) # (!\Mux21~1_combout  & (\Mux85~3_combout  & !\Add0~19 )))

	.dataa(Mux21),
	.datab(Mux85),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~19 ),
	.combout(\Add0~20_combout ),
	.cout(\Add0~21 ));
// synopsys translate_off
defparam \Add0~20 .lut_mask = 16'h698E;
defparam \Add0~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N6
cycloneive_lcell_comb \aluif.portOut[10]~106 (
// Equation(s):
// \aluif.portOut[10]~106_combout  = (\aluif.portOut[10]~105_combout  & ((\prif.ALUOP_ex [1]) # ((\portOut~30_combout )))) # (!\aluif.portOut[10]~105_combout  & (!\prif.ALUOP_ex [1] & ((\Add0~20_combout ))))

	.dataa(\aluif.portOut[10]~105_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\portOut~30_combout ),
	.datad(\Add0~20_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[10]~106_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[10]~106 .lut_mask = 16'hB9A8;
defparam \aluif.portOut[10]~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N4
cycloneive_lcell_comb \aluif.portOut[10]~107 (
// Equation(s):
// \aluif.portOut[10]~107_combout  = (\aluif.portOut[15]~80_combout  & ((\Add1~20_combout ) # ((\aluif.portOut[15]~86_combout )))) # (!\aluif.portOut[15]~80_combout  & (((!\aluif.portOut[15]~86_combout  & \aluif.portOut[10]~106_combout ))))

	.dataa(\Add1~20_combout ),
	.datab(\aluif.portOut[15]~80_combout ),
	.datac(\aluif.portOut[15]~86_combout ),
	.datad(\aluif.portOut[10]~106_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[10]~107_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[10]~107 .lut_mask = 16'hCBC8;
defparam \aluif.portOut[10]~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N0
cycloneive_lcell_comb \ShiftRight0~108 (
// Equation(s):
// \ShiftRight0~108_combout  = (!\Mux92~2_combout  & ((\Mux93~2_combout  & ((\ShiftRight0~77_combout ))) # (!\Mux93~2_combout  & (\ShiftRight0~79_combout ))))

	.dataa(\ShiftRight0~79_combout ),
	.datab(Mux92),
	.datac(Mux931),
	.datad(\ShiftRight0~77_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~108_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~108 .lut_mask = 16'h3202;
defparam \ShiftRight0~108 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N16
cycloneive_lcell_comb \aluif.portOut[10]~103 (
// Equation(s):
// \aluif.portOut[10]~103_combout  = (\aluif.portOut[15]~82_combout  & ((\aluif.portOut[15]~83_combout  & (\portOut~29_combout )) # (!\aluif.portOut[15]~83_combout  & ((\ShiftRight0~108_combout ))))) # (!\aluif.portOut[15]~82_combout  & 
// (((\aluif.portOut[15]~83_combout ))))

	.dataa(\portOut~29_combout ),
	.datab(\ShiftRight0~108_combout ),
	.datac(\aluif.portOut[15]~82_combout ),
	.datad(\aluif.portOut[15]~83_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[10]~103_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[10]~103 .lut_mask = 16'hAFC0;
defparam \aluif.portOut[10]~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N10
cycloneive_lcell_comb \aluif.portOut[10]~104 (
// Equation(s):
// \aluif.portOut[10]~104_combout  = (\aluif.portOut[10]~103_combout  & (((\aluif.portOut[15]~81_combout ) # (\ShiftRight0~85_combout )))) # (!\aluif.portOut[10]~103_combout  & (\ShiftRight0~91_combout  & (!\aluif.portOut[15]~81_combout )))

	.dataa(\ShiftRight0~91_combout ),
	.datab(\aluif.portOut[10]~103_combout ),
	.datac(\aluif.portOut[15]~81_combout ),
	.datad(\ShiftRight0~85_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[10]~104_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[10]~104 .lut_mask = 16'hCEC2;
defparam \aluif.portOut[10]~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N4
cycloneive_lcell_comb \ShiftRight0~109 (
// Equation(s):
// \ShiftRight0~109_combout  = (\ShiftRight0~61_combout  & ((\ShiftRight0~26_combout ) # ((\Mux2~1_combout  & \ShiftLeft0~16_combout ))))

	.dataa(Mux2),
	.datab(\ShiftLeft0~16_combout ),
	.datac(\ShiftRight0~61_combout ),
	.datad(\ShiftRight0~26_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~109_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~109 .lut_mask = 16'hF080;
defparam \ShiftRight0~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y23_N4
cycloneive_lcell_comb \portOut~32 (
// Equation(s):
// \portOut~32_combout  = (\Mux18~1_combout ) # (\Mux82~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux18),
	.datad(Mux82),
	.cin(gnd),
	.combout(\portOut~32_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~32 .lut_mask = 16'hFFF0;
defparam \portOut~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N18
cycloneive_lcell_comb \aluif.portOut[13]~109 (
// Equation(s):
// \aluif.portOut[13]~109_combout  = (\aluif.portOut[15]~83_combout  & (((\portOut~32_combout )) # (!\aluif.portOut[15]~82_combout ))) # (!\aluif.portOut[15]~83_combout  & (\aluif.portOut[15]~82_combout  & (\ShiftRight0~109_combout )))

	.dataa(\aluif.portOut[15]~83_combout ),
	.datab(\aluif.portOut[15]~82_combout ),
	.datac(\ShiftRight0~109_combout ),
	.datad(\portOut~32_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[13]~109_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[13]~109 .lut_mask = 16'hEA62;
defparam \aluif.portOut[13]~109 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N12
cycloneive_lcell_comb \aluif.portOut[13]~110 (
// Equation(s):
// \aluif.portOut[13]~110_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[13]~109_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[13]~109_combout  & (\ShiftRight0~94_combout )) # (!\aluif.portOut[13]~109_combout  & 
// ((\ShiftRight0~92_combout )))))

	.dataa(\ShiftRight0~94_combout ),
	.datab(\aluif.portOut[15]~81_combout ),
	.datac(\ShiftRight0~92_combout ),
	.datad(\aluif.portOut[13]~109_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[13]~110_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[13]~110 .lut_mask = 16'hEE30;
defparam \aluif.portOut[13]~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y23_N6
cycloneive_lcell_comb \portOut~33 (
// Equation(s):
// \portOut~33_combout  = \Mux18~1_combout  $ (\Mux82~3_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux18),
	.datad(Mux82),
	.cin(gnd),
	.combout(\portOut~33_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~33 .lut_mask = 16'h0FF0;
defparam \portOut~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y22_N4
cycloneive_lcell_comb \ShiftLeft0~53 (
// Equation(s):
// \ShiftLeft0~53_combout  = (\Mux92~2_combout  & ((\Mux93~2_combout  & ((\ShiftLeft0~22_combout ))) # (!\Mux93~2_combout  & (\ShiftLeft0~24_combout ))))

	.dataa(Mux931),
	.datab(Mux92),
	.datac(\ShiftLeft0~24_combout ),
	.datad(\ShiftLeft0~22_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~53_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~53 .lut_mask = 16'hC840;
defparam \ShiftLeft0~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N26
cycloneive_lcell_comb \ShiftLeft0~45 (
// Equation(s):
// \ShiftLeft0~45_combout  = (\Mux95~1_combout  & ((\Mux21~1_combout ))) # (!\Mux95~1_combout  & (\Mux20~1_combout ))

	.dataa(gnd),
	.datab(Mux95),
	.datac(Mux20),
	.datad(Mux21),
	.cin(gnd),
	.combout(\ShiftLeft0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~45 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N6
cycloneive_lcell_comb \ShiftLeft0~55 (
// Equation(s):
// \ShiftLeft0~55_combout  = (\Mux94~1_combout  & ((\ShiftLeft0~45_combout ))) # (!\Mux94~1_combout  & (\ShiftLeft0~54_combout ))

	.dataa(\ShiftLeft0~54_combout ),
	.datab(gnd),
	.datac(\ShiftLeft0~45_combout ),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftLeft0~55_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~55 .lut_mask = 16'hF0AA;
defparam \ShiftLeft0~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N6
cycloneive_lcell_comb \ShiftLeft0~56 (
// Equation(s):
// \ShiftLeft0~56_combout  = (\Mux93~2_combout  & (\ShiftLeft0~38_combout )) # (!\Mux93~2_combout  & ((\ShiftLeft0~55_combout )))

	.dataa(Mux931),
	.datab(gnd),
	.datac(\ShiftLeft0~38_combout ),
	.datad(\ShiftLeft0~55_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~56_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~56 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N28
cycloneive_lcell_comb \ShiftLeft0~57 (
// Equation(s):
// \ShiftLeft0~57_combout  = (\ShiftLeft0~53_combout ) # ((!\Mux92~2_combout  & \ShiftLeft0~56_combout ))

	.dataa(Mux92),
	.datab(gnd),
	.datac(\ShiftLeft0~53_combout ),
	.datad(\ShiftLeft0~56_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~57_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~57 .lut_mask = 16'hF5F0;
defparam \ShiftLeft0~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N12
cycloneive_lcell_comb \aluif.portOut[13]~111 (
// Equation(s):
// \aluif.portOut[13]~111_combout  = (\prif.ALUOP_ex [2] & (((\ShiftLeft0~57_combout  & \aluif.portOut[15]~26_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~34_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(\portOut~34_combout ),
	.datab(\ShiftLeft0~57_combout ),
	.datac(prifALUOP_ex_2),
	.datad(\aluif.portOut[15]~26_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[13]~111_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[13]~111 .lut_mask = 16'hCA0F;
defparam \aluif.portOut[13]~111 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N26
cycloneive_lcell_comb \aluif.portOut[13]~112 (
// Equation(s):
// \aluif.portOut[13]~112_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[13]~111_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[13]~111_combout  & ((\portOut~33_combout ))) # (!\aluif.portOut[13]~111_combout  & (\Add0~26_combout ))))

	.dataa(\Add0~26_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\portOut~33_combout ),
	.datad(\aluif.portOut[13]~111_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[13]~112_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[13]~112 .lut_mask = 16'hFC22;
defparam \aluif.portOut[13]~112 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N24
cycloneive_lcell_comb \Add1~24 (
// Equation(s):
// \Add1~24_combout  = ((\Mux19~3_combout  $ (\Mux83~3_combout  $ (\Add1~23 )))) # (GND)
// \Add1~25  = CARRY((\Mux19~3_combout  & ((!\Add1~23 ) # (!\Mux83~3_combout ))) # (!\Mux19~3_combout  & (!\Mux83~3_combout  & !\Add1~23 )))

	.dataa(Mux192),
	.datab(Mux83),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~23 ),
	.combout(\Add1~24_combout ),
	.cout(\Add1~25 ));
// synopsys translate_off
defparam \Add1~24 .lut_mask = 16'h962B;
defparam \Add1~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N26
cycloneive_lcell_comb \Add1~26 (
// Equation(s):
// \Add1~26_combout  = (\Mux82~3_combout  & ((\Mux18~1_combout  & (!\Add1~25 )) # (!\Mux18~1_combout  & ((\Add1~25 ) # (GND))))) # (!\Mux82~3_combout  & ((\Mux18~1_combout  & (\Add1~25  & VCC)) # (!\Mux18~1_combout  & (!\Add1~25 ))))
// \Add1~27  = CARRY((\Mux82~3_combout  & ((!\Add1~25 ) # (!\Mux18~1_combout ))) # (!\Mux82~3_combout  & (!\Mux18~1_combout  & !\Add1~25 )))

	.dataa(Mux82),
	.datab(Mux18),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~25 ),
	.combout(\Add1~26_combout ),
	.cout(\Add1~27 ));
// synopsys translate_off
defparam \Add1~26 .lut_mask = 16'h692B;
defparam \Add1~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N20
cycloneive_lcell_comb \aluif.portOut[13]~113 (
// Equation(s):
// \aluif.portOut[13]~113_combout  = (\aluif.portOut[15]~80_combout  & (((\aluif.portOut[15]~86_combout ) # (\Add1~26_combout )))) # (!\aluif.portOut[15]~80_combout  & (\aluif.portOut[13]~112_combout  & (!\aluif.portOut[15]~86_combout )))

	.dataa(\aluif.portOut[13]~112_combout ),
	.datab(\aluif.portOut[15]~80_combout ),
	.datac(\aluif.portOut[15]~86_combout ),
	.datad(\Add1~26_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[13]~113_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[13]~113 .lut_mask = 16'hCEC2;
defparam \aluif.portOut[13]~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N8
cycloneive_lcell_comb \portOut~35 (
// Equation(s):
// \portOut~35_combout  = (\Mux19~0_combout ) # ((\Mux83~3_combout ) # (\Mux19~1_combout ))

	.dataa(Mux19),
	.datab(gnd),
	.datac(Mux83),
	.datad(Mux191),
	.cin(gnd),
	.combout(\portOut~35_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~35 .lut_mask = 16'hFFFA;
defparam \portOut~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N24
cycloneive_lcell_comb \Add0~24 (
// Equation(s):
// \Add0~24_combout  = ((\Mux83~3_combout  $ (\Mux19~3_combout  $ (!\Add0~23 )))) # (GND)
// \Add0~25  = CARRY((\Mux83~3_combout  & ((\Mux19~3_combout ) # (!\Add0~23 ))) # (!\Mux83~3_combout  & (\Mux19~3_combout  & !\Add0~23 )))

	.dataa(Mux83),
	.datab(Mux192),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~23 ),
	.combout(\Add0~24_combout ),
	.cout(\Add0~25 ));
// synopsys translate_off
defparam \Add0~24 .lut_mask = 16'h698E;
defparam \Add0~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N16
cycloneive_lcell_comb \ShiftLeft0~58 (
// Equation(s):
// \ShiftLeft0~58_combout  = (\Mux93~2_combout  & (\Mux31~1_combout  & (\ShiftLeft0~16_combout ))) # (!\Mux93~2_combout  & (((\ShiftLeft0~28_combout ))))

	.dataa(Mux31),
	.datab(\ShiftLeft0~16_combout ),
	.datac(\ShiftLeft0~28_combout ),
	.datad(Mux931),
	.cin(gnd),
	.combout(\ShiftLeft0~58_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~58 .lut_mask = 16'h88F0;
defparam \ShiftLeft0~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y23_N24
cycloneive_lcell_comb \ShiftLeft0~62 (
// Equation(s):
// \ShiftLeft0~62_combout  = (\Mux92~2_combout  & ((\ShiftLeft0~58_combout ))) # (!\Mux92~2_combout  & (\ShiftLeft0~61_combout ))

	.dataa(\ShiftLeft0~61_combout ),
	.datab(gnd),
	.datac(Mux92),
	.datad(\ShiftLeft0~58_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~62_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~62 .lut_mask = 16'hFA0A;
defparam \ShiftLeft0~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N8
cycloneive_lcell_comb \aluif.portOut[12]~117 (
// Equation(s):
// \aluif.portOut[12]~117_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[15]~26_combout  & \ShiftLeft0~62_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~37_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(\portOut~37_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\ShiftLeft0~62_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[12]~117_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[12]~117 .lut_mask = 16'hE323;
defparam \aluif.portOut[12]~117 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N12
cycloneive_lcell_comb \portOut~36 (
// Equation(s):
// \portOut~36_combout  = \Mux83~3_combout  $ (((\Mux19~1_combout ) # (\Mux19~0_combout )))

	.dataa(Mux191),
	.datab(gnd),
	.datac(Mux83),
	.datad(Mux19),
	.cin(gnd),
	.combout(\portOut~36_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~36 .lut_mask = 16'h0F5A;
defparam \portOut~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N14
cycloneive_lcell_comb \aluif.portOut[12]~118 (
// Equation(s):
// \aluif.portOut[12]~118_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[12]~117_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[12]~117_combout  & ((\portOut~36_combout ))) # (!\aluif.portOut[12]~117_combout  & (\Add0~24_combout ))))

	.dataa(prifALUOP_ex_1),
	.datab(\Add0~24_combout ),
	.datac(\aluif.portOut[12]~117_combout ),
	.datad(\portOut~36_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[12]~118_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[12]~118 .lut_mask = 16'hF4A4;
defparam \aluif.portOut[12]~118 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N28
cycloneive_lcell_comb \ShiftRight0~39 (
// Equation(s):
// \ShiftRight0~39_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux4~1_combout )) # (!\Mux95~1_combout  & ((\Mux5~1_combout ))))) # (!\Mux94~1_combout  & (((\Mux95~1_combout ))))

	.dataa(Mux4),
	.datab(Mux5),
	.datac(Mux94),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftRight0~39_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~39 .lut_mask = 16'hAFC0;
defparam \ShiftRight0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N14
cycloneive_lcell_comb \ShiftRight0~40 (
// Equation(s):
// \ShiftRight0~40_combout  = (\Mux94~1_combout  & (((\ShiftRight0~39_combout )))) # (!\Mux94~1_combout  & ((\ShiftRight0~39_combout  & ((\Mux6~1_combout ))) # (!\ShiftRight0~39_combout  & (\Mux7~1_combout ))))

	.dataa(Mux7),
	.datab(Mux94),
	.datac(Mux6),
	.datad(\ShiftRight0~39_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~40_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~40 .lut_mask = 16'hFC22;
defparam \ShiftRight0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N12
cycloneive_lcell_comb \ShiftRight0~97 (
// Equation(s):
// \ShiftRight0~97_combout  = (\Mux93~2_combout  & (((\ShiftRight0~40_combout )))) # (!\Mux93~2_combout  & ((\ShiftRight0~37_combout ) # ((\ShiftRight0~36_combout ))))

	.dataa(\ShiftRight0~37_combout ),
	.datab(\ShiftRight0~36_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~40_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~97 .lut_mask = 16'hFE0E;
defparam \ShiftRight0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N4
cycloneive_lcell_comb \ShiftRight0~42 (
// Equation(s):
// \ShiftRight0~42_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux2~1_combout ))) # (!\Mux95~1_combout  & (\Mux3~1_combout ))))

	.dataa(Mux3),
	.datab(Mux95),
	.datac(Mux2),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftRight0~42_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~42 .lut_mask = 16'h00E2;
defparam \ShiftRight0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N8
cycloneive_lcell_comb \ShiftRight0~110 (
// Equation(s):
// \ShiftRight0~110_combout  = (\ShiftRight0~61_combout  & ((\ShiftRight0~42_combout ) # ((\Mux94~1_combout  & \ShiftRight0~43_combout ))))

	.dataa(Mux94),
	.datab(\ShiftRight0~61_combout ),
	.datac(\ShiftRight0~42_combout ),
	.datad(\ShiftRight0~43_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~110_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~110 .lut_mask = 16'hC8C0;
defparam \ShiftRight0~110 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N24
cycloneive_lcell_comb \aluif.portOut[12]~115 (
// Equation(s):
// \aluif.portOut[12]~115_combout  = (\aluif.portOut[15]~82_combout  & ((\aluif.portOut[15]~83_combout  & (\portOut~35_combout )) # (!\aluif.portOut[15]~83_combout  & ((\ShiftRight0~110_combout ))))) # (!\aluif.portOut[15]~82_combout  & 
// (((\aluif.portOut[15]~83_combout ))))

	.dataa(\portOut~35_combout ),
	.datab(\ShiftRight0~110_combout ),
	.datac(\aluif.portOut[15]~82_combout ),
	.datad(\aluif.portOut[15]~83_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[12]~115_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[12]~115 .lut_mask = 16'hAFC0;
defparam \aluif.portOut[12]~115 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N2
cycloneive_lcell_comb \aluif.portOut[12]~116 (
// Equation(s):
// \aluif.portOut[12]~116_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[12]~115_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[12]~115_combout  & ((\ShiftRight0~97_combout ))) # (!\aluif.portOut[12]~115_combout  & 
// (\ShiftRight0~96_combout ))))

	.dataa(\ShiftRight0~96_combout ),
	.datab(\aluif.portOut[15]~81_combout ),
	.datac(\ShiftRight0~97_combout ),
	.datad(\aluif.portOut[12]~115_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[12]~116_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[12]~116 .lut_mask = 16'hFC22;
defparam \aluif.portOut[12]~116 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N16
cycloneive_lcell_comb \aluif.portOut[12]~119 (
// Equation(s):
// \aluif.portOut[12]~119_combout  = (\aluif.portOut[15]~86_combout  & (((\aluif.portOut[15]~80_combout ) # (\aluif.portOut[12]~116_combout )))) # (!\aluif.portOut[15]~86_combout  & (\aluif.portOut[12]~118_combout  & (!\aluif.portOut[15]~80_combout )))

	.dataa(\aluif.portOut[15]~86_combout ),
	.datab(\aluif.portOut[12]~118_combout ),
	.datac(\aluif.portOut[15]~80_combout ),
	.datad(\aluif.portOut[12]~116_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[12]~119_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[12]~119 .lut_mask = 16'hAEA4;
defparam \aluif.portOut[12]~119 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N22
cycloneive_lcell_comb \portOut~38 (
// Equation(s):
// \portOut~38_combout  = (\Mux80~4_combout ) # (\Mux16~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux80),
	.datad(Mux16),
	.cin(gnd),
	.combout(\portOut~38_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~38 .lut_mask = 16'hFFF0;
defparam \portOut~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N28
cycloneive_lcell_comb \Add1~28 (
// Equation(s):
// \Add1~28_combout  = ((\Mux81~3_combout  $ (\Mux17~1_combout  $ (\Add1~27 )))) # (GND)
// \Add1~29  = CARRY((\Mux81~3_combout  & (\Mux17~1_combout  & !\Add1~27 )) # (!\Mux81~3_combout  & ((\Mux17~1_combout ) # (!\Add1~27 ))))

	.dataa(Mux81),
	.datab(Mux17),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~27 ),
	.combout(\Add1~28_combout ),
	.cout(\Add1~29 ));
// synopsys translate_off
defparam \Add1~28 .lut_mask = 16'h964D;
defparam \Add1~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y25_N30
cycloneive_lcell_comb \Add1~30 (
// Equation(s):
// \Add1~30_combout  = (\Mux16~1_combout  & ((\Mux80~4_combout  & (!\Add1~29 )) # (!\Mux80~4_combout  & (\Add1~29  & VCC)))) # (!\Mux16~1_combout  & ((\Mux80~4_combout  & ((\Add1~29 ) # (GND))) # (!\Mux80~4_combout  & (!\Add1~29 ))))
// \Add1~31  = CARRY((\Mux16~1_combout  & (\Mux80~4_combout  & !\Add1~29 )) # (!\Mux16~1_combout  & ((\Mux80~4_combout ) # (!\Add1~29 ))))

	.dataa(Mux16),
	.datab(Mux80),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~29 ),
	.combout(\Add1~30_combout ),
	.cout(\Add1~31 ));
// synopsys translate_off
defparam \Add1~30 .lut_mask = 16'h694D;
defparam \Add1~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N28
cycloneive_lcell_comb \portOut~39 (
// Equation(s):
// \portOut~39_combout  = \Mux80~4_combout  $ (\Mux16~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux80),
	.datad(Mux16),
	.cin(gnd),
	.combout(\portOut~39_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~39 .lut_mask = 16'h0FF0;
defparam \portOut~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N28
cycloneive_lcell_comb \Add0~28 (
// Equation(s):
// \Add0~28_combout  = ((\Mux17~1_combout  $ (\Mux81~3_combout  $ (!\Add0~27 )))) # (GND)
// \Add0~29  = CARRY((\Mux17~1_combout  & ((\Mux81~3_combout ) # (!\Add0~27 ))) # (!\Mux17~1_combout  & (\Mux81~3_combout  & !\Add0~27 )))

	.dataa(Mux17),
	.datab(Mux81),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~27 ),
	.combout(\Add0~28_combout ),
	.cout(\Add0~29 ));
// synopsys translate_off
defparam \Add0~28 .lut_mask = 16'h698E;
defparam \Add0~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y25_N30
cycloneive_lcell_comb \Add0~30 (
// Equation(s):
// \Add0~30_combout  = (\Mux16~1_combout  & ((\Mux80~4_combout  & (\Add0~29  & VCC)) # (!\Mux80~4_combout  & (!\Add0~29 )))) # (!\Mux16~1_combout  & ((\Mux80~4_combout  & (!\Add0~29 )) # (!\Mux80~4_combout  & ((\Add0~29 ) # (GND)))))
// \Add0~31  = CARRY((\Mux16~1_combout  & (!\Mux80~4_combout  & !\Add0~29 )) # (!\Mux16~1_combout  & ((!\Add0~29 ) # (!\Mux80~4_combout ))))

	.dataa(Mux16),
	.datab(Mux80),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~29 ),
	.combout(\Add0~30_combout ),
	.cout(\Add0~31 ));
// synopsys translate_off
defparam \Add0~30 .lut_mask = 16'h9617;
defparam \Add0~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N16
cycloneive_lcell_comb \ShiftLeft0~63 (
// Equation(s):
// \ShiftLeft0~63_combout  = (\Mux92~2_combout  & ((\Mux93~2_combout  & ((\ShiftLeft0~30_combout ))) # (!\Mux93~2_combout  & (\ShiftLeft0~32_combout ))))

	.dataa(\ShiftLeft0~32_combout ),
	.datab(Mux92),
	.datac(Mux931),
	.datad(\ShiftLeft0~30_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~63_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~63 .lut_mask = 16'hC808;
defparam \ShiftLeft0~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N10
cycloneive_lcell_comb \ShiftLeft0~54 (
// Equation(s):
// \ShiftLeft0~54_combout  = (\Mux95~1_combout  & ((\Mux19~1_combout ) # ((\Mux19~0_combout )))) # (!\Mux95~1_combout  & (((\Mux18~1_combout ))))

	.dataa(Mux191),
	.datab(Mux95),
	.datac(Mux18),
	.datad(Mux19),
	.cin(gnd),
	.combout(\ShiftLeft0~54_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~54 .lut_mask = 16'hFCB8;
defparam \ShiftLeft0~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N6
cycloneive_lcell_comb \ShiftLeft0~64 (
// Equation(s):
// \ShiftLeft0~64_combout  = (\Mux95~1_combout  & ((\Mux17~1_combout ))) # (!\Mux95~1_combout  & (\Mux16~1_combout ))

	.dataa(Mux95),
	.datab(gnd),
	.datac(Mux16),
	.datad(Mux17),
	.cin(gnd),
	.combout(\ShiftLeft0~64_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~64 .lut_mask = 16'hFA50;
defparam \ShiftLeft0~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N24
cycloneive_lcell_comb \ShiftLeft0~65 (
// Equation(s):
// \ShiftLeft0~65_combout  = (\Mux94~1_combout  & (\ShiftLeft0~54_combout )) # (!\Mux94~1_combout  & ((\ShiftLeft0~64_combout )))

	.dataa(Mux94),
	.datab(gnd),
	.datac(\ShiftLeft0~54_combout ),
	.datad(\ShiftLeft0~64_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~65_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~65 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N2
cycloneive_lcell_comb \ShiftLeft0~66 (
// Equation(s):
// \ShiftLeft0~66_combout  = (\Mux93~2_combout  & ((\ShiftLeft0~46_combout ))) # (!\Mux93~2_combout  & (\ShiftLeft0~65_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~65_combout ),
	.datac(\ShiftLeft0~46_combout ),
	.datad(Mux931),
	.cin(gnd),
	.combout(\ShiftLeft0~66_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~66 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N12
cycloneive_lcell_comb \ShiftLeft0~67 (
// Equation(s):
// \ShiftLeft0~67_combout  = (\ShiftLeft0~63_combout ) # ((!\Mux92~2_combout  & \ShiftLeft0~66_combout ))

	.dataa(gnd),
	.datab(Mux92),
	.datac(\ShiftLeft0~63_combout ),
	.datad(\ShiftLeft0~66_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~67_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~67 .lut_mask = 16'hF3F0;
defparam \ShiftLeft0~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N10
cycloneive_lcell_comb \portOut~40 (
// Equation(s):
// \portOut~40_combout  = (\Mux80~4_combout  & \Mux16~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux80),
	.datad(Mux16),
	.cin(gnd),
	.combout(\portOut~40_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~40 .lut_mask = 16'hF000;
defparam \portOut~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N24
cycloneive_lcell_comb \aluif.portOut[15]~123 (
// Equation(s):
// \aluif.portOut[15]~123_combout  = (\prif.ALUOP_ex [2] & (\aluif.portOut[15]~26_combout  & (\ShiftLeft0~67_combout ))) # (!\prif.ALUOP_ex [2] & (((\portOut~40_combout )) # (!\aluif.portOut[15]~26_combout )))

	.dataa(prifALUOP_ex_2),
	.datab(\aluif.portOut[15]~26_combout ),
	.datac(\ShiftLeft0~67_combout ),
	.datad(\portOut~40_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[15]~123_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~123 .lut_mask = 16'hD591;
defparam \aluif.portOut[15]~123 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N18
cycloneive_lcell_comb \aluif.portOut[15]~124 (
// Equation(s):
// \aluif.portOut[15]~124_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[15]~123_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[15]~123_combout  & (\portOut~39_combout )) # (!\aluif.portOut[15]~123_combout  & ((\Add0~30_combout )))))

	.dataa(prifALUOP_ex_1),
	.datab(\portOut~39_combout ),
	.datac(\Add0~30_combout ),
	.datad(\aluif.portOut[15]~123_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[15]~124_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~124 .lut_mask = 16'hEE50;
defparam \aluif.portOut[15]~124 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N8
cycloneive_lcell_comb \aluif.portOut[15]~125 (
// Equation(s):
// \aluif.portOut[15]~125_combout  = (\aluif.portOut[15]~80_combout  & ((\aluif.portOut[15]~86_combout ) # ((\Add1~30_combout )))) # (!\aluif.portOut[15]~80_combout  & (!\aluif.portOut[15]~86_combout  & ((\aluif.portOut[15]~124_combout ))))

	.dataa(\aluif.portOut[15]~80_combout ),
	.datab(\aluif.portOut[15]~86_combout ),
	.datac(\Add1~30_combout ),
	.datad(\aluif.portOut[15]~124_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[15]~125_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~125 .lut_mask = 16'hB9A8;
defparam \aluif.portOut[15]~125 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N18
cycloneive_lcell_comb \ShiftRight0~113 (
// Equation(s):
// \ShiftRight0~113_combout  = (!\Mux94~1_combout  & (!\Mux95~1_combout  & (\Mux0~1_combout  & \ShiftRight0~61_combout )))

	.dataa(Mux94),
	.datab(Mux95),
	.datac(Mux0),
	.datad(\ShiftRight0~61_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~113_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~113 .lut_mask = 16'h1000;
defparam \ShiftRight0~113 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N12
cycloneive_lcell_comb \aluif.portOut[15]~121 (
// Equation(s):
// \aluif.portOut[15]~121_combout  = (\aluif.portOut[15]~83_combout  & ((\portOut~38_combout ) # ((!\aluif.portOut[15]~82_combout )))) # (!\aluif.portOut[15]~83_combout  & (((\ShiftRight0~113_combout  & \aluif.portOut[15]~82_combout ))))

	.dataa(\portOut~38_combout ),
	.datab(\aluif.portOut[15]~83_combout ),
	.datac(\ShiftRight0~113_combout ),
	.datad(\aluif.portOut[15]~82_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[15]~121_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~121 .lut_mask = 16'hB8CC;
defparam \aluif.portOut[15]~121 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y24_N2
cycloneive_lcell_comb \aluif.portOut[15]~122 (
// Equation(s):
// \aluif.portOut[15]~122_combout  = (\aluif.portOut[15]~121_combout  & ((\aluif.portOut[15]~81_combout ) # ((\ShiftRight0~100_combout )))) # (!\aluif.portOut[15]~121_combout  & (!\aluif.portOut[15]~81_combout  & (\ShiftRight0~99_combout )))

	.dataa(\aluif.portOut[15]~121_combout ),
	.datab(\aluif.portOut[15]~81_combout ),
	.datac(\ShiftRight0~99_combout ),
	.datad(\ShiftRight0~100_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[15]~122_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[15]~122 .lut_mask = 16'hBA98;
defparam \aluif.portOut[15]~122 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N30
cycloneive_lcell_comb \portOut~41 (
// Equation(s):
// \portOut~41_combout  = (\Mux81~3_combout ) # (\Mux17~1_combout )

	.dataa(Mux81),
	.datab(gnd),
	.datac(Mux17),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~41_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~41 .lut_mask = 16'hFAFA;
defparam \portOut~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N4
cycloneive_lcell_comb \portOut~43 (
// Equation(s):
// \portOut~43_combout  = (\Mux81~3_combout  & \Mux17~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux81),
	.datad(Mux17),
	.cin(gnd),
	.combout(\portOut~43_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~43 .lut_mask = 16'hF000;
defparam \portOut~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N6
cycloneive_lcell_comb \aluif.portOut[14]~129 (
// Equation(s):
// \aluif.portOut[14]~129_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & (\ShiftLeft0~72_combout )) # (!\prif.ALUOP_ex [2] & ((\portOut~43_combout ))))) # (!\aluif.portOut[15]~26_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\ShiftLeft0~72_combout ),
	.datab(\portOut~43_combout ),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(prifALUOP_ex_2),
	.cin(gnd),
	.combout(\aluif.portOut[14]~129_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[14]~129 .lut_mask = 16'hA0CF;
defparam \aluif.portOut[14]~129 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N20
cycloneive_lcell_comb \aluif.portOut[14]~130 (
// Equation(s):
// \aluif.portOut[14]~130_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[14]~129_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[14]~129_combout  & (\portOut~42_combout )) # (!\aluif.portOut[14]~129_combout  & ((\Add0~28_combout )))))

	.dataa(\portOut~42_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\Add0~28_combout ),
	.datad(\aluif.portOut[14]~129_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[14]~130_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[14]~130 .lut_mask = 16'hEE30;
defparam \aluif.portOut[14]~130 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N28
cycloneive_lcell_comb \aluif.portOut[14]~128 (
// Equation(s):
// \aluif.portOut[14]~128_combout  = (\aluif.portOut[14]~127_combout  & (((\ShiftRight0~103_combout ) # (\aluif.portOut[15]~81_combout )))) # (!\aluif.portOut[14]~127_combout  & (\ShiftRight0~102_combout  & ((!\aluif.portOut[15]~81_combout ))))

	.dataa(\aluif.portOut[14]~127_combout ),
	.datab(\ShiftRight0~102_combout ),
	.datac(\ShiftRight0~103_combout ),
	.datad(\aluif.portOut[15]~81_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[14]~128_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[14]~128 .lut_mask = 16'hAAE4;
defparam \aluif.portOut[14]~128 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N2
cycloneive_lcell_comb \aluif.portOut[14]~131 (
// Equation(s):
// \aluif.portOut[14]~131_combout  = (\aluif.portOut[15]~80_combout  & (((\aluif.portOut[15]~86_combout )))) # (!\aluif.portOut[15]~80_combout  & ((\aluif.portOut[15]~86_combout  & ((\aluif.portOut[14]~128_combout ))) # (!\aluif.portOut[15]~86_combout  & 
// (\aluif.portOut[14]~130_combout ))))

	.dataa(\aluif.portOut[14]~130_combout ),
	.datab(\aluif.portOut[15]~80_combout ),
	.datac(\aluif.portOut[15]~86_combout ),
	.datad(\aluif.portOut[14]~128_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[14]~131_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[14]~131 .lut_mask = 16'hF2C2;
defparam \aluif.portOut[14]~131 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N0
cycloneive_lcell_comb \Add1~32 (
// Equation(s):
// \Add1~32_combout  = ((\Mux79~0_combout  $ (\Mux15~1_combout  $ (\Add1~31 )))) # (GND)
// \Add1~33  = CARRY((\Mux79~0_combout  & (\Mux15~1_combout  & !\Add1~31 )) # (!\Mux79~0_combout  & ((\Mux15~1_combout ) # (!\Add1~31 ))))

	.dataa(Mux79),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~31 ),
	.combout(\Add1~32_combout ),
	.cout(\Add1~33 ));
// synopsys translate_off
defparam \Add1~32 .lut_mask = 16'h964D;
defparam \Add1~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N2
cycloneive_lcell_comb \Add1~34 (
// Equation(s):
// \Add1~34_combout  = (\Mux78~0_combout  & ((\Mux14~1_combout  & (!\Add1~33 )) # (!\Mux14~1_combout  & ((\Add1~33 ) # (GND))))) # (!\Mux78~0_combout  & ((\Mux14~1_combout  & (\Add1~33  & VCC)) # (!\Mux14~1_combout  & (!\Add1~33 ))))
// \Add1~35  = CARRY((\Mux78~0_combout  & ((!\Add1~33 ) # (!\Mux14~1_combout ))) # (!\Mux78~0_combout  & (!\Mux14~1_combout  & !\Add1~33 )))

	.dataa(Mux78),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~33 ),
	.combout(\Add1~34_combout ),
	.cout(\Add1~35 ));
// synopsys translate_off
defparam \Add1~34 .lut_mask = 16'h692B;
defparam \Add1~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N4
cycloneive_lcell_comb \Add1~36 (
// Equation(s):
// \Add1~36_combout  = ((\Mux77~0_combout  $ (\Mux13~1_combout  $ (\Add1~35 )))) # (GND)
// \Add1~37  = CARRY((\Mux77~0_combout  & (\Mux13~1_combout  & !\Add1~35 )) # (!\Mux77~0_combout  & ((\Mux13~1_combout ) # (!\Add1~35 ))))

	.dataa(Mux77),
	.datab(Mux13),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~35 ),
	.combout(\Add1~36_combout ),
	.cout(\Add1~37 ));
// synopsys translate_off
defparam \Add1~36 .lut_mask = 16'h964D;
defparam \Add1~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N6
cycloneive_lcell_comb \Add1~38 (
// Equation(s):
// \Add1~38_combout  = (\Mux76~0_combout  & ((\Mux12~1_combout  & (!\Add1~37 )) # (!\Mux12~1_combout  & ((\Add1~37 ) # (GND))))) # (!\Mux76~0_combout  & ((\Mux12~1_combout  & (\Add1~37  & VCC)) # (!\Mux12~1_combout  & (!\Add1~37 ))))
// \Add1~39  = CARRY((\Mux76~0_combout  & ((!\Add1~37 ) # (!\Mux12~1_combout ))) # (!\Mux76~0_combout  & (!\Mux12~1_combout  & !\Add1~37 )))

	.dataa(Mux76),
	.datab(Mux12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~37 ),
	.combout(\Add1~38_combout ),
	.cout(\Add1~39 ));
// synopsys translate_off
defparam \Add1~38 .lut_mask = 16'h692B;
defparam \Add1~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N8
cycloneive_lcell_comb \Add1~40 (
// Equation(s):
// \Add1~40_combout  = ((\Mux11~1_combout  $ (\Mux75~0_combout  $ (\Add1~39 )))) # (GND)
// \Add1~41  = CARRY((\Mux11~1_combout  & ((!\Add1~39 ) # (!\Mux75~0_combout ))) # (!\Mux11~1_combout  & (!\Mux75~0_combout  & !\Add1~39 )))

	.dataa(Mux11),
	.datab(Mux75),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~39 ),
	.combout(\Add1~40_combout ),
	.cout(\Add1~41 ));
// synopsys translate_off
defparam \Add1~40 .lut_mask = 16'h962B;
defparam \Add1~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N10
cycloneive_lcell_comb \Add1~42 (
// Equation(s):
// \Add1~42_combout  = (\Mux74~0_combout  & ((\Mux10~1_combout  & (!\Add1~41 )) # (!\Mux10~1_combout  & ((\Add1~41 ) # (GND))))) # (!\Mux74~0_combout  & ((\Mux10~1_combout  & (\Add1~41  & VCC)) # (!\Mux10~1_combout  & (!\Add1~41 ))))
// \Add1~43  = CARRY((\Mux74~0_combout  & ((!\Add1~41 ) # (!\Mux10~1_combout ))) # (!\Mux74~0_combout  & (!\Mux10~1_combout  & !\Add1~41 )))

	.dataa(Mux74),
	.datab(Mux10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~41 ),
	.combout(\Add1~42_combout ),
	.cout(\Add1~43 ));
// synopsys translate_off
defparam \Add1~42 .lut_mask = 16'h692B;
defparam \Add1~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N12
cycloneive_lcell_comb \Add1~44 (
// Equation(s):
// \Add1~44_combout  = ((\Mux73~0_combout  $ (\Mux9~1_combout  $ (\Add1~43 )))) # (GND)
// \Add1~45  = CARRY((\Mux73~0_combout  & (\Mux9~1_combout  & !\Add1~43 )) # (!\Mux73~0_combout  & ((\Mux9~1_combout ) # (!\Add1~43 ))))

	.dataa(Mux73),
	.datab(Mux9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~43 ),
	.combout(\Add1~44_combout ),
	.cout(\Add1~45 ));
// synopsys translate_off
defparam \Add1~44 .lut_mask = 16'h964D;
defparam \Add1~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N14
cycloneive_lcell_comb \Add1~46 (
// Equation(s):
// \Add1~46_combout  = (\Mux8~1_combout  & ((\Mux72~0_combout  & (!\Add1~45 )) # (!\Mux72~0_combout  & (\Add1~45  & VCC)))) # (!\Mux8~1_combout  & ((\Mux72~0_combout  & ((\Add1~45 ) # (GND))) # (!\Mux72~0_combout  & (!\Add1~45 ))))
// \Add1~47  = CARRY((\Mux8~1_combout  & (\Mux72~0_combout  & !\Add1~45 )) # (!\Mux8~1_combout  & ((\Mux72~0_combout ) # (!\Add1~45 ))))

	.dataa(Mux8),
	.datab(Mux72),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~45 ),
	.combout(\Add1~46_combout ),
	.cout(\Add1~47 ));
// synopsys translate_off
defparam \Add1~46 .lut_mask = 16'h694D;
defparam \Add1~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N18
cycloneive_lcell_comb \portOut~44 (
// Equation(s):
// \portOut~44_combout  = (\Mux8~1_combout ) # (\Mux72~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux8),
	.datad(Mux72),
	.cin(gnd),
	.combout(\portOut~44_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~44 .lut_mask = 16'hFFF0;
defparam \portOut~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N16
cycloneive_lcell_comb \aluif.portOut[23]~133 (
// Equation(s):
// \aluif.portOut[23]~133_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & (\ShiftRight0~101_combout )) # (!\prif.ALUOP_ex [2] & ((\portOut~44_combout ))))) # (!\aluif.portOut[15]~26_combout  & (!\prif.ALUOP_ex [2]))

	.dataa(\aluif.portOut[15]~26_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\ShiftRight0~101_combout ),
	.datad(\portOut~44_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[23]~133_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[23]~133 .lut_mask = 16'hB391;
defparam \aluif.portOut[23]~133 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N26
cycloneive_lcell_comb \aluif.portOut[23]~134 (
// Equation(s):
// \aluif.portOut[23]~134_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[23]~133_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[23]~133_combout  & ((!\portOut~44_combout ))) # (!\aluif.portOut[23]~133_combout  & (\Add1~46_combout ))))

	.dataa(\Add1~46_combout ),
	.datab(\portOut~44_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.portOut[23]~133_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[23]~134_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[23]~134 .lut_mask = 16'hF30A;
defparam \aluif.portOut[23]~134 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N0
cycloneive_lcell_comb \portOut~46 (
// Equation(s):
// \portOut~46_combout  = \Mux8~1_combout  $ (\Mux72~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux8),
	.datad(Mux72),
	.cin(gnd),
	.combout(\portOut~46_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~46 .lut_mask = 16'h0FF0;
defparam \portOut~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N10
cycloneive_lcell_comb \aluif.portOut[23]~135 (
// Equation(s):
// \aluif.portOut[23]~135_combout  = ((!\prif.ALUOP_ex [2] & !\prif.ALUOP_ex [1])) # (!\prif.ALUOP_ex [0])

	.dataa(prifALUOP_ex_0),
	.datab(prifALUOP_ex_2),
	.datac(prifALUOP_ex_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\aluif.portOut[23]~135_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[23]~135 .lut_mask = 16'h5757;
defparam \aluif.portOut[23]~135 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N28
cycloneive_lcell_comb \aluif.portOut[23]~136 (
// Equation(s):
// \aluif.portOut[23]~136_combout  = (!\prif.ALUOP_ex [1] & \prif.ALUOP_ex [0])

	.dataa(gnd),
	.datab(gnd),
	.datac(prifALUOP_ex_1),
	.datad(prifALUOP_ex_0),
	.cin(gnd),
	.combout(\aluif.portOut[23]~136_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[23]~136 .lut_mask = 16'h0F00;
defparam \aluif.portOut[23]~136 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N0
cycloneive_lcell_comb \ShiftLeft0~75 (
// Equation(s):
// \ShiftLeft0~75_combout  = (\Mux95~1_combout  & ((\Mux94~1_combout  & ((\Mux15~1_combout ))) # (!\Mux94~1_combout  & (\Mux13~1_combout ))))

	.dataa(Mux94),
	.datab(Mux13),
	.datac(Mux95),
	.datad(Mux15),
	.cin(gnd),
	.combout(\ShiftLeft0~75_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~75 .lut_mask = 16'hE040;
defparam \ShiftLeft0~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N2
cycloneive_lcell_comb \ShiftLeft0~73 (
// Equation(s):
// \ShiftLeft0~73_combout  = (\Mux95~1_combout  & (((\Mux94~1_combout )))) # (!\Mux95~1_combout  & ((\Mux94~1_combout  & (\Mux10~1_combout )) # (!\Mux94~1_combout  & ((\Mux8~1_combout )))))

	.dataa(Mux95),
	.datab(Mux10),
	.datac(Mux8),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftLeft0~73_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~73 .lut_mask = 16'hEE50;
defparam \ShiftLeft0~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N0
cycloneive_lcell_comb \ShiftLeft0~74 (
// Equation(s):
// \ShiftLeft0~74_combout  = (\Mux95~1_combout  & ((\ShiftLeft0~73_combout  & ((\Mux11~1_combout ))) # (!\ShiftLeft0~73_combout  & (\Mux9~1_combout )))) # (!\Mux95~1_combout  & (((\ShiftLeft0~73_combout ))))

	.dataa(Mux9),
	.datab(Mux95),
	.datac(Mux11),
	.datad(\ShiftLeft0~73_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~74_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~74 .lut_mask = 16'hF388;
defparam \ShiftLeft0~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N18
cycloneive_lcell_comb \ShiftLeft0~77 (
// Equation(s):
// \ShiftLeft0~77_combout  = (\Mux93~2_combout  & ((\ShiftLeft0~76_combout ) # ((\ShiftLeft0~75_combout )))) # (!\Mux93~2_combout  & (((\ShiftLeft0~74_combout ))))

	.dataa(\ShiftLeft0~76_combout ),
	.datab(Mux931),
	.datac(\ShiftLeft0~75_combout ),
	.datad(\ShiftLeft0~74_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~77_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~77 .lut_mask = 16'hFBC8;
defparam \ShiftLeft0~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N4
cycloneive_lcell_comb \portOut~45 (
// Equation(s):
// \portOut~45_combout  = (\Mux8~1_combout  & \Mux72~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux8),
	.datad(Mux72),
	.cin(gnd),
	.combout(\portOut~45_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~45 .lut_mask = 16'hF000;
defparam \portOut~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N2
cycloneive_lcell_comb \aluif.portOut[23]~137 (
// Equation(s):
// \aluif.portOut[23]~137_combout  = (\aluif.portOut[15]~83_combout  & ((\portOut~45_combout ) # ((!\aluif.portOut[15]~82_combout )))) # (!\aluif.portOut[15]~83_combout  & (((\aluif.portOut[15]~82_combout  & \ShiftLeft0~33_combout ))))

	.dataa(\aluif.portOut[15]~83_combout ),
	.datab(\portOut~45_combout ),
	.datac(\aluif.portOut[15]~82_combout ),
	.datad(\ShiftLeft0~33_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[23]~137_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[23]~137 .lut_mask = 16'hDA8A;
defparam \aluif.portOut[23]~137 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N8
cycloneive_lcell_comb \aluif.portOut[23]~138 (
// Equation(s):
// \aluif.portOut[23]~138_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[23]~137_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[23]~137_combout  & (\ShiftLeft0~66_combout )) # (!\aluif.portOut[23]~137_combout  & 
// ((\ShiftLeft0~77_combout )))))

	.dataa(\ShiftLeft0~66_combout ),
	.datab(\aluif.portOut[15]~81_combout ),
	.datac(\ShiftLeft0~77_combout ),
	.datad(\aluif.portOut[23]~137_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[23]~138_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[23]~138 .lut_mask = 16'hEE30;
defparam \aluif.portOut[23]~138 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N0
cycloneive_lcell_comb \Add0~32 (
// Equation(s):
// \Add0~32_combout  = ((\Mux79~0_combout  $ (\Mux15~1_combout  $ (!\Add0~31 )))) # (GND)
// \Add0~33  = CARRY((\Mux79~0_combout  & ((\Mux15~1_combout ) # (!\Add0~31 ))) # (!\Mux79~0_combout  & (\Mux15~1_combout  & !\Add0~31 )))

	.dataa(Mux79),
	.datab(Mux15),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~31 ),
	.combout(\Add0~32_combout ),
	.cout(\Add0~33 ));
// synopsys translate_off
defparam \Add0~32 .lut_mask = 16'h698E;
defparam \Add0~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N2
cycloneive_lcell_comb \Add0~34 (
// Equation(s):
// \Add0~34_combout  = (\Mux78~0_combout  & ((\Mux14~1_combout  & (\Add0~33  & VCC)) # (!\Mux14~1_combout  & (!\Add0~33 )))) # (!\Mux78~0_combout  & ((\Mux14~1_combout  & (!\Add0~33 )) # (!\Mux14~1_combout  & ((\Add0~33 ) # (GND)))))
// \Add0~35  = CARRY((\Mux78~0_combout  & (!\Mux14~1_combout  & !\Add0~33 )) # (!\Mux78~0_combout  & ((!\Add0~33 ) # (!\Mux14~1_combout ))))

	.dataa(Mux78),
	.datab(Mux14),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~33 ),
	.combout(\Add0~34_combout ),
	.cout(\Add0~35 ));
// synopsys translate_off
defparam \Add0~34 .lut_mask = 16'h9617;
defparam \Add0~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N4
cycloneive_lcell_comb \Add0~36 (
// Equation(s):
// \Add0~36_combout  = ((\Mux13~1_combout  $ (\Mux77~0_combout  $ (!\Add0~35 )))) # (GND)
// \Add0~37  = CARRY((\Mux13~1_combout  & ((\Mux77~0_combout ) # (!\Add0~35 ))) # (!\Mux13~1_combout  & (\Mux77~0_combout  & !\Add0~35 )))

	.dataa(Mux13),
	.datab(Mux77),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~35 ),
	.combout(\Add0~36_combout ),
	.cout(\Add0~37 ));
// synopsys translate_off
defparam \Add0~36 .lut_mask = 16'h698E;
defparam \Add0~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N6
cycloneive_lcell_comb \Add0~38 (
// Equation(s):
// \Add0~38_combout  = (\Mux76~0_combout  & ((\Mux12~1_combout  & (\Add0~37  & VCC)) # (!\Mux12~1_combout  & (!\Add0~37 )))) # (!\Mux76~0_combout  & ((\Mux12~1_combout  & (!\Add0~37 )) # (!\Mux12~1_combout  & ((\Add0~37 ) # (GND)))))
// \Add0~39  = CARRY((\Mux76~0_combout  & (!\Mux12~1_combout  & !\Add0~37 )) # (!\Mux76~0_combout  & ((!\Add0~37 ) # (!\Mux12~1_combout ))))

	.dataa(Mux76),
	.datab(Mux12),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~37 ),
	.combout(\Add0~38_combout ),
	.cout(\Add0~39 ));
// synopsys translate_off
defparam \Add0~38 .lut_mask = 16'h9617;
defparam \Add0~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N8
cycloneive_lcell_comb \Add0~40 (
// Equation(s):
// \Add0~40_combout  = ((\Mux11~1_combout  $ (\Mux75~0_combout  $ (!\Add0~39 )))) # (GND)
// \Add0~41  = CARRY((\Mux11~1_combout  & ((\Mux75~0_combout ) # (!\Add0~39 ))) # (!\Mux11~1_combout  & (\Mux75~0_combout  & !\Add0~39 )))

	.dataa(Mux11),
	.datab(Mux75),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~39 ),
	.combout(\Add0~40_combout ),
	.cout(\Add0~41 ));
// synopsys translate_off
defparam \Add0~40 .lut_mask = 16'h698E;
defparam \Add0~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N10
cycloneive_lcell_comb \Add0~42 (
// Equation(s):
// \Add0~42_combout  = (\Mux74~0_combout  & ((\Mux10~1_combout  & (\Add0~41  & VCC)) # (!\Mux10~1_combout  & (!\Add0~41 )))) # (!\Mux74~0_combout  & ((\Mux10~1_combout  & (!\Add0~41 )) # (!\Mux10~1_combout  & ((\Add0~41 ) # (GND)))))
// \Add0~43  = CARRY((\Mux74~0_combout  & (!\Mux10~1_combout  & !\Add0~41 )) # (!\Mux74~0_combout  & ((!\Add0~41 ) # (!\Mux10~1_combout ))))

	.dataa(Mux74),
	.datab(Mux10),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~41 ),
	.combout(\Add0~42_combout ),
	.cout(\Add0~43 ));
// synopsys translate_off
defparam \Add0~42 .lut_mask = 16'h9617;
defparam \Add0~42 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N12
cycloneive_lcell_comb \Add0~44 (
// Equation(s):
// \Add0~44_combout  = ((\Mux73~0_combout  $ (\Mux9~1_combout  $ (!\Add0~43 )))) # (GND)
// \Add0~45  = CARRY((\Mux73~0_combout  & ((\Mux9~1_combout ) # (!\Add0~43 ))) # (!\Mux73~0_combout  & (\Mux9~1_combout  & !\Add0~43 )))

	.dataa(Mux73),
	.datab(Mux9),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~43 ),
	.combout(\Add0~44_combout ),
	.cout(\Add0~45 ));
// synopsys translate_off
defparam \Add0~44 .lut_mask = 16'h698E;
defparam \Add0~44 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N14
cycloneive_lcell_comb \Add0~46 (
// Equation(s):
// \Add0~46_combout  = (\Mux72~0_combout  & ((\Mux8~1_combout  & (\Add0~45  & VCC)) # (!\Mux8~1_combout  & (!\Add0~45 )))) # (!\Mux72~0_combout  & ((\Mux8~1_combout  & (!\Add0~45 )) # (!\Mux8~1_combout  & ((\Add0~45 ) # (GND)))))
// \Add0~47  = CARRY((\Mux72~0_combout  & (!\Mux8~1_combout  & !\Add0~45 )) # (!\Mux72~0_combout  & ((!\Add0~45 ) # (!\Mux8~1_combout ))))

	.dataa(Mux72),
	.datab(Mux8),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~45 ),
	.combout(\Add0~46_combout ),
	.cout(\Add0~47 ));
// synopsys translate_off
defparam \Add0~46 .lut_mask = 16'h9617;
defparam \Add0~46 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N6
cycloneive_lcell_comb \aluif.portOut[23]~139 (
// Equation(s):
// \aluif.portOut[23]~139_combout  = (\aluif.portOut[23]~136_combout  & ((\aluif.portOut[23]~135_combout ) # ((\Add0~46_combout )))) # (!\aluif.portOut[23]~136_combout  & (!\aluif.portOut[23]~135_combout  & (\aluif.portOut[23]~138_combout )))

	.dataa(\aluif.portOut[23]~136_combout ),
	.datab(\aluif.portOut[23]~135_combout ),
	.datac(\aluif.portOut[23]~138_combout ),
	.datad(\Add0~46_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[23]~139_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[23]~139 .lut_mask = 16'hBA98;
defparam \aluif.portOut[23]~139 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N30
cycloneive_lcell_comb \aluif.portOut[22]~144 (
// Equation(s):
// \aluif.portOut[22]~144_combout  = (\aluif.portOut[23]~135_combout  & ((\Mux73~0_combout  $ (!\Mux9~1_combout )) # (!\aluif.portOut[23]~136_combout )))

	.dataa(\aluif.portOut[23]~135_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(Mux73),
	.datad(Mux9),
	.cin(gnd),
	.combout(\aluif.portOut[22]~144_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~144 .lut_mask = 16'hA22A;
defparam \aluif.portOut[22]~144 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N2
cycloneive_lcell_comb \portOut~48 (
// Equation(s):
// \portOut~48_combout  = (\Mux73~0_combout ) # (\Mux9~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux73),
	.datad(Mux9),
	.cin(gnd),
	.combout(\portOut~48_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~48 .lut_mask = 16'hFFF0;
defparam \portOut~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N20
cycloneive_lcell_comb \aluif.portOut[22]~143 (
// Equation(s):
// \aluif.portOut[22]~143_combout  = (\prif.ALUOP_ex [2] & (\aluif.portOut[15]~26_combout  & (\ShiftRight0~104_combout ))) # (!\prif.ALUOP_ex [2] & (((\portOut~48_combout )) # (!\aluif.portOut[15]~26_combout )))

	.dataa(prifALUOP_ex_2),
	.datab(\aluif.portOut[15]~26_combout ),
	.datac(\ShiftRight0~104_combout ),
	.datad(\portOut~48_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[22]~143_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~143 .lut_mask = 16'hD591;
defparam \aluif.portOut[22]~143 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N26
cycloneive_lcell_comb \aluif.portOut[22]~259 (
// Equation(s):
// \aluif.portOut[22]~259_combout  = (\aluif.portOut[22]~143_combout  & ((\prif.ALUOP_ex [1]) # ((!\Mux9~1_combout  & !\Mux73~0_combout ))))

	.dataa(Mux9),
	.datab(prifALUOP_ex_1),
	.datac(Mux73),
	.datad(\aluif.portOut[22]~143_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[22]~259_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~259 .lut_mask = 16'hCD00;
defparam \aluif.portOut[22]~259 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N24
cycloneive_lcell_comb \ShiftLeft0~49 (
// Equation(s):
// \ShiftLeft0~49_combout  = (\Mux95~1_combout  & (\Mux22~1_combout )) # (!\Mux95~1_combout  & ((\Mux21~1_combout )))

	.dataa(Mux95),
	.datab(gnd),
	.datac(Mux22),
	.datad(Mux21),
	.cin(gnd),
	.combout(\ShiftLeft0~49_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~49 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N28
cycloneive_lcell_comb \ShiftLeft0~50 (
// Equation(s):
// \ShiftLeft0~50_combout  = (\Mux94~1_combout  & (\ShiftLeft0~41_combout )) # (!\Mux94~1_combout  & ((\ShiftLeft0~49_combout )))

	.dataa(Mux94),
	.datab(gnd),
	.datac(\ShiftLeft0~41_combout ),
	.datad(\ShiftLeft0~49_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~50_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~50 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y24_N18
cycloneive_lcell_comb \ShiftLeft0~59 (
// Equation(s):
// \ShiftLeft0~59_combout  = (\Mux95~1_combout  & (((\Mux20~1_combout )))) # (!\Mux95~1_combout  & ((\Mux19~1_combout ) # ((\Mux19~0_combout ))))

	.dataa(Mux191),
	.datab(Mux95),
	.datac(Mux20),
	.datad(Mux19),
	.cin(gnd),
	.combout(\ShiftLeft0~59_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~59 .lut_mask = 16'hF3E2;
defparam \ShiftLeft0~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N12
cycloneive_lcell_comb \ShiftLeft0~69 (
// Equation(s):
// \ShiftLeft0~69_combout  = (\Mux95~1_combout  & ((\Mux18~1_combout ))) # (!\Mux95~1_combout  & (\Mux17~1_combout ))

	.dataa(gnd),
	.datab(Mux95),
	.datac(Mux17),
	.datad(Mux18),
	.cin(gnd),
	.combout(\ShiftLeft0~69_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~69 .lut_mask = 16'hFC30;
defparam \ShiftLeft0~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N6
cycloneive_lcell_comb \ShiftLeft0~70 (
// Equation(s):
// \ShiftLeft0~70_combout  = (\Mux94~1_combout  & (\ShiftLeft0~59_combout )) # (!\Mux94~1_combout  & ((\ShiftLeft0~69_combout )))

	.dataa(Mux94),
	.datab(gnd),
	.datac(\ShiftLeft0~59_combout ),
	.datad(\ShiftLeft0~69_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~70_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~70 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N20
cycloneive_lcell_comb \ShiftLeft0~71 (
// Equation(s):
// \ShiftLeft0~71_combout  = (\Mux93~2_combout  & (\ShiftLeft0~50_combout )) # (!\Mux93~2_combout  & ((\ShiftLeft0~70_combout )))

	.dataa(gnd),
	.datab(\ShiftLeft0~50_combout ),
	.datac(Mux931),
	.datad(\ShiftLeft0~70_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~71_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~71 .lut_mask = 16'hCFC0;
defparam \ShiftLeft0~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N8
cycloneive_lcell_comb \portOut~47 (
// Equation(s):
// \portOut~47_combout  = (\Mux73~0_combout  & \Mux9~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux73),
	.datad(Mux9),
	.cin(gnd),
	.combout(\portOut~47_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~47 .lut_mask = 16'hF000;
defparam \portOut~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N14
cycloneive_lcell_comb \aluif.portOut[22]~141 (
// Equation(s):
// \aluif.portOut[22]~141_combout  = (\aluif.portOut[15]~82_combout  & ((\aluif.portOut[15]~83_combout  & ((\portOut~47_combout ))) # (!\aluif.portOut[15]~83_combout  & (\ShiftLeft0~36_combout )))) # (!\aluif.portOut[15]~82_combout  & 
// (((\aluif.portOut[15]~83_combout ))))

	.dataa(\ShiftLeft0~36_combout ),
	.datab(\portOut~47_combout ),
	.datac(\aluif.portOut[15]~82_combout ),
	.datad(\aluif.portOut[15]~83_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[22]~141_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~141 .lut_mask = 16'hCFA0;
defparam \aluif.portOut[22]~141 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N4
cycloneive_lcell_comb \ShiftLeft0~80 (
// Equation(s):
// \ShiftLeft0~80_combout  = (\Mux95~1_combout  & ((\Mux94~1_combout  & (\Mux16~1_combout )) # (!\Mux94~1_combout  & ((\Mux14~1_combout )))))

	.dataa(Mux16),
	.datab(Mux14),
	.datac(Mux95),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftLeft0~80_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~80 .lut_mask = 16'hA0C0;
defparam \ShiftLeft0~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N14
cycloneive_lcell_comb \ShiftLeft0~79 (
// Equation(s):
// \ShiftLeft0~79_combout  = (\ShiftLeft0~78_combout  & (((\Mux12~1_combout ) # (!\Mux95~1_combout )))) # (!\ShiftLeft0~78_combout  & (\Mux10~1_combout  & (\Mux95~1_combout )))

	.dataa(\ShiftLeft0~78_combout ),
	.datab(Mux10),
	.datac(Mux95),
	.datad(Mux12),
	.cin(gnd),
	.combout(\ShiftLeft0~79_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~79 .lut_mask = 16'hEA4A;
defparam \ShiftLeft0~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N2
cycloneive_lcell_comb \ShiftLeft0~81 (
// Equation(s):
// \ShiftLeft0~81_combout  = (!\Mux95~1_combout  & ((\Mux94~1_combout  & ((\Mux15~1_combout ))) # (!\Mux94~1_combout  & (\Mux13~1_combout ))))

	.dataa(Mux94),
	.datab(Mux13),
	.datac(Mux95),
	.datad(Mux15),
	.cin(gnd),
	.combout(\ShiftLeft0~81_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~81 .lut_mask = 16'h0E04;
defparam \ShiftLeft0~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N16
cycloneive_lcell_comb \ShiftLeft0~82 (
// Equation(s):
// \ShiftLeft0~82_combout  = (\Mux93~2_combout  & ((\ShiftLeft0~80_combout ) # ((\ShiftLeft0~81_combout )))) # (!\Mux93~2_combout  & (((\ShiftLeft0~79_combout ))))

	.dataa(Mux931),
	.datab(\ShiftLeft0~80_combout ),
	.datac(\ShiftLeft0~79_combout ),
	.datad(\ShiftLeft0~81_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~82_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~82 .lut_mask = 16'hFAD8;
defparam \ShiftLeft0~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N16
cycloneive_lcell_comb \aluif.portOut[22]~142 (
// Equation(s):
// \aluif.portOut[22]~142_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[22]~141_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[22]~141_combout  & (\ShiftLeft0~71_combout )) # (!\aluif.portOut[22]~141_combout  & 
// ((\ShiftLeft0~82_combout )))))

	.dataa(\aluif.portOut[15]~81_combout ),
	.datab(\ShiftLeft0~71_combout ),
	.datac(\aluif.portOut[22]~141_combout ),
	.datad(\ShiftLeft0~82_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[22]~142_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~142 .lut_mask = 16'hE5E0;
defparam \aluif.portOut[22]~142 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N12
cycloneive_lcell_comb \aluif.portOut[22]~145 (
// Equation(s):
// \aluif.portOut[22]~145_combout  = (\aluif.portOut[22]~144_combout  & (!\aluif.portOut[23]~136_combout  & (\aluif.portOut[22]~259_combout ))) # (!\aluif.portOut[22]~144_combout  & ((\aluif.portOut[23]~136_combout ) # ((\aluif.portOut[22]~142_combout ))))

	.dataa(\aluif.portOut[22]~144_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(\aluif.portOut[22]~259_combout ),
	.datad(\aluif.portOut[22]~142_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[22]~145_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~145 .lut_mask = 16'h7564;
defparam \aluif.portOut[22]~145 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N4
cycloneive_lcell_comb \aluif.portOut[22]~260 (
// Equation(s):
// \aluif.portOut[22]~260_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[22]~143_combout )))) # (!\prif.ALUOP_ex [1] & (((!\Mux9~1_combout  & !\Mux73~0_combout )) # (!\aluif.portOut[22]~143_combout )))

	.dataa(Mux9),
	.datab(prifALUOP_ex_1),
	.datac(Mux73),
	.datad(\aluif.portOut[22]~143_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[22]~260_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~260 .lut_mask = 16'hCD33;
defparam \aluif.portOut[22]~260 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N18
cycloneive_lcell_comb \aluif.portOut[22]~146 (
// Equation(s):
// \aluif.portOut[22]~146_combout  = (\aluif.portOut[23]~135_combout  & (!\aluif.portOut[23]~136_combout  & (\aluif.portOut[22]~260_combout ))) # (!\aluif.portOut[23]~135_combout  & ((\aluif.portOut[23]~136_combout ) # ((\aluif.portOut[22]~142_combout ))))

	.dataa(\aluif.portOut[23]~135_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(\aluif.portOut[22]~260_combout ),
	.datad(\aluif.portOut[22]~142_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[22]~146_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~146 .lut_mask = 16'h7564;
defparam \aluif.portOut[22]~146 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N6
cycloneive_lcell_comb \aluif.portOut[22]~261 (
// Equation(s):
// \aluif.portOut[22]~261_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[22]~146_combout )))) # (!\prif.ALUOP_ex [1] & ((\prif.ALUOP_ex [0] & (\aluif.portOut[22]~145_combout  & !\aluif.portOut[22]~146_combout )) # (!\prif.ALUOP_ex [0] & 
// ((\aluif.portOut[22]~146_combout )))))

	.dataa(\aluif.portOut[22]~145_combout ),
	.datab(prifALUOP_ex_1),
	.datac(prifALUOP_ex_0),
	.datad(\aluif.portOut[22]~146_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[22]~261_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[22]~261 .lut_mask = 16'hCF20;
defparam \aluif.portOut[22]~261 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N2
cycloneive_lcell_comb \portOut~51 (
// Equation(s):
// \portOut~51_combout  = \Mux74~0_combout  $ (\Mux10~1_combout )

	.dataa(gnd),
	.datab(Mux74),
	.datac(gnd),
	.datad(Mux10),
	.cin(gnd),
	.combout(\portOut~51_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~51 .lut_mask = 16'h33CC;
defparam \portOut~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N30
cycloneive_lcell_comb \portOut~49 (
// Equation(s):
// \portOut~49_combout  = (\Mux10~1_combout ) # (\Mux74~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux10),
	.datad(Mux74),
	.cin(gnd),
	.combout(\portOut~49_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~49 .lut_mask = 16'hFFF0;
defparam \portOut~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N20
cycloneive_lcell_comb \aluif.portOut[21]~148 (
// Equation(s):
// \aluif.portOut[21]~148_combout  = (\prif.ALUOP_ex [2] & (\ShiftRight0~95_combout  & ((\aluif.portOut[15]~26_combout )))) # (!\prif.ALUOP_ex [2] & (((\portOut~49_combout ) # (!\aluif.portOut[15]~26_combout ))))

	.dataa(\ShiftRight0~95_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\portOut~49_combout ),
	.datad(\aluif.portOut[15]~26_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[21]~148_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[21]~148 .lut_mask = 16'hB833;
defparam \aluif.portOut[21]~148 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N22
cycloneive_lcell_comb \aluif.portOut[21]~149 (
// Equation(s):
// \aluif.portOut[21]~149_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[21]~148_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[21]~148_combout  & (!\portOut~49_combout )) # (!\aluif.portOut[21]~148_combout  & ((\Add1~42_combout )))))

	.dataa(\portOut~49_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\Add1~42_combout ),
	.datad(\aluif.portOut[21]~148_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[21]~149_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[21]~149 .lut_mask = 16'hDD30;
defparam \aluif.portOut[21]~149 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N30
cycloneive_lcell_comb \ShiftLeft0~83 (
// Equation(s):
// \ShiftLeft0~83_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux15~1_combout )) # (!\Mux95~1_combout  & ((\Mux14~1_combout )))))

	.dataa(Mux15),
	.datab(Mux94),
	.datac(Mux14),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftLeft0~83_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~83 .lut_mask = 16'h2230;
defparam \ShiftLeft0~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N24
cycloneive_lcell_comb \ShiftLeft0~84 (
// Equation(s):
// \ShiftLeft0~84_combout  = (\ShiftLeft0~83_combout ) # ((\Mux94~1_combout  & \ShiftLeft0~64_combout ))

	.dataa(gnd),
	.datab(Mux94),
	.datac(\ShiftLeft0~83_combout ),
	.datad(\ShiftLeft0~64_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~84_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~84 .lut_mask = 16'hFCF0;
defparam \ShiftLeft0~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N18
cycloneive_lcell_comb \ShiftLeft0~85 (
// Equation(s):
// \ShiftLeft0~85_combout  = (\Mux95~1_combout  & (\Mux94~1_combout )) # (!\Mux95~1_combout  & ((\Mux94~1_combout  & ((\Mux12~1_combout ))) # (!\Mux94~1_combout  & (\Mux10~1_combout ))))

	.dataa(Mux95),
	.datab(Mux94),
	.datac(Mux10),
	.datad(Mux12),
	.cin(gnd),
	.combout(\ShiftLeft0~85_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~85 .lut_mask = 16'hDC98;
defparam \ShiftLeft0~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N20
cycloneive_lcell_comb \ShiftLeft0~86 (
// Equation(s):
// \ShiftLeft0~86_combout  = (\Mux95~1_combout  & ((\ShiftLeft0~85_combout  & ((\Mux13~1_combout ))) # (!\ShiftLeft0~85_combout  & (\Mux11~1_combout )))) # (!\Mux95~1_combout  & (((\ShiftLeft0~85_combout ))))

	.dataa(Mux11),
	.datab(Mux13),
	.datac(Mux95),
	.datad(\ShiftLeft0~85_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~86_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~86 .lut_mask = 16'hCFA0;
defparam \ShiftLeft0~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N16
cycloneive_lcell_comb \ShiftLeft0~87 (
// Equation(s):
// \ShiftLeft0~87_combout  = (\Mux93~2_combout  & (\ShiftLeft0~84_combout )) # (!\Mux93~2_combout  & ((\ShiftLeft0~86_combout )))

	.dataa(Mux931),
	.datab(gnd),
	.datac(\ShiftLeft0~84_combout ),
	.datad(\ShiftLeft0~86_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~87_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~87 .lut_mask = 16'hF5A0;
defparam \ShiftLeft0~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N18
cycloneive_lcell_comb \portOut~50 (
// Equation(s):
// \portOut~50_combout  = (\Mux10~1_combout  & \Mux74~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux10),
	.datad(Mux74),
	.cin(gnd),
	.combout(\portOut~50_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~50 .lut_mask = 16'hF000;
defparam \portOut~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N4
cycloneive_lcell_comb \aluif.portOut[21]~150 (
// Equation(s):
// \aluif.portOut[21]~150_combout  = (\aluif.portOut[15]~83_combout  & ((\portOut~50_combout ) # ((!\aluif.portOut[15]~82_combout )))) # (!\aluif.portOut[15]~83_combout  & (((\aluif.portOut[15]~82_combout  & \ShiftLeft0~25_combout ))))

	.dataa(\aluif.portOut[15]~83_combout ),
	.datab(\portOut~50_combout ),
	.datac(\aluif.portOut[15]~82_combout ),
	.datad(\ShiftLeft0~25_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[21]~150_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[21]~150 .lut_mask = 16'hDA8A;
defparam \aluif.portOut[21]~150 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N2
cycloneive_lcell_comb \aluif.portOut[21]~151 (
// Equation(s):
// \aluif.portOut[21]~151_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[21]~150_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[21]~150_combout  & ((\ShiftLeft0~56_combout ))) # (!\aluif.portOut[21]~150_combout  & 
// (\ShiftLeft0~87_combout ))))

	.dataa(\aluif.portOut[15]~81_combout ),
	.datab(\ShiftLeft0~87_combout ),
	.datac(\aluif.portOut[21]~150_combout ),
	.datad(\ShiftLeft0~56_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[21]~151_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[21]~151 .lut_mask = 16'hF4A4;
defparam \aluif.portOut[21]~151 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N24
cycloneive_lcell_comb \aluif.portOut[21]~152 (
// Equation(s):
// \aluif.portOut[21]~152_combout  = (\aluif.portOut[23]~136_combout  & ((\aluif.portOut[23]~135_combout ) # ((\Add0~42_combout )))) # (!\aluif.portOut[23]~136_combout  & (!\aluif.portOut[23]~135_combout  & ((\aluif.portOut[21]~151_combout ))))

	.dataa(\aluif.portOut[23]~136_combout ),
	.datab(\aluif.portOut[23]~135_combout ),
	.datac(\Add0~42_combout ),
	.datad(\aluif.portOut[21]~151_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[21]~152_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[21]~152 .lut_mask = 16'hB9A8;
defparam \aluif.portOut[21]~152 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N26
cycloneive_lcell_comb \aluif.portOut[28]~154 (
// Equation(s):
// \aluif.portOut[28]~154_combout  = (\aluif.portOut[5]~25_combout  & (!\aluif.portOut[2]~32_combout  & ((!\ShiftLeft0~15_combout ) # (!\aluif.portOut[1]~13_combout ))))

	.dataa(\aluif.portOut[1]~13_combout ),
	.datab(\aluif.portOut[5]~25_combout ),
	.datac(\ShiftLeft0~15_combout ),
	.datad(\aluif.portOut[2]~32_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~154_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~154 .lut_mask = 16'h004C;
defparam \aluif.portOut[28]~154 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N16
cycloneive_lcell_comb \Add1~48 (
// Equation(s):
// \Add1~48_combout  = ((\Mux7~1_combout  $ (\Mux71~0_combout  $ (\Add1~47 )))) # (GND)
// \Add1~49  = CARRY((\Mux7~1_combout  & ((!\Add1~47 ) # (!\Mux71~0_combout ))) # (!\Mux7~1_combout  & (!\Mux71~0_combout  & !\Add1~47 )))

	.dataa(Mux7),
	.datab(Mux71),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~47 ),
	.combout(\Add1~48_combout ),
	.cout(\Add1~49 ));
// synopsys translate_off
defparam \Add1~48 .lut_mask = 16'h962B;
defparam \Add1~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N18
cycloneive_lcell_comb \Add1~50 (
// Equation(s):
// \Add1~50_combout  = (\Mux70~0_combout  & ((\Mux6~1_combout  & (!\Add1~49 )) # (!\Mux6~1_combout  & ((\Add1~49 ) # (GND))))) # (!\Mux70~0_combout  & ((\Mux6~1_combout  & (\Add1~49  & VCC)) # (!\Mux6~1_combout  & (!\Add1~49 ))))
// \Add1~51  = CARRY((\Mux70~0_combout  & ((!\Add1~49 ) # (!\Mux6~1_combout ))) # (!\Mux70~0_combout  & (!\Mux6~1_combout  & !\Add1~49 )))

	.dataa(Mux70),
	.datab(Mux6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~49 ),
	.combout(\Add1~50_combout ),
	.cout(\Add1~51 ));
// synopsys translate_off
defparam \Add1~50 .lut_mask = 16'h692B;
defparam \Add1~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N20
cycloneive_lcell_comb \Add1~52 (
// Equation(s):
// \Add1~52_combout  = ((\Mux5~1_combout  $ (\Mux69~0_combout  $ (\Add1~51 )))) # (GND)
// \Add1~53  = CARRY((\Mux5~1_combout  & ((!\Add1~51 ) # (!\Mux69~0_combout ))) # (!\Mux5~1_combout  & (!\Mux69~0_combout  & !\Add1~51 )))

	.dataa(Mux5),
	.datab(Mux69),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~51 ),
	.combout(\Add1~52_combout ),
	.cout(\Add1~53 ));
// synopsys translate_off
defparam \Add1~52 .lut_mask = 16'h962B;
defparam \Add1~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N22
cycloneive_lcell_comb \Add1~54 (
// Equation(s):
// \Add1~54_combout  = (\Mux68~0_combout  & ((\Mux4~1_combout  & (!\Add1~53 )) # (!\Mux4~1_combout  & ((\Add1~53 ) # (GND))))) # (!\Mux68~0_combout  & ((\Mux4~1_combout  & (\Add1~53  & VCC)) # (!\Mux4~1_combout  & (!\Add1~53 ))))
// \Add1~55  = CARRY((\Mux68~0_combout  & ((!\Add1~53 ) # (!\Mux4~1_combout ))) # (!\Mux68~0_combout  & (!\Mux4~1_combout  & !\Add1~53 )))

	.dataa(Mux68),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~53 ),
	.combout(\Add1~54_combout ),
	.cout(\Add1~55 ));
// synopsys translate_off
defparam \Add1~54 .lut_mask = 16'h692B;
defparam \Add1~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N24
cycloneive_lcell_comb \Add1~56 (
// Equation(s):
// \Add1~56_combout  = ((\Mux3~1_combout  $ (\Mux67~0_combout  $ (\Add1~55 )))) # (GND)
// \Add1~57  = CARRY((\Mux3~1_combout  & ((!\Add1~55 ) # (!\Mux67~0_combout ))) # (!\Mux3~1_combout  & (!\Mux67~0_combout  & !\Add1~55 )))

	.dataa(Mux3),
	.datab(Mux67),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~55 ),
	.combout(\Add1~56_combout ),
	.cout(\Add1~57 ));
// synopsys translate_off
defparam \Add1~56 .lut_mask = 16'h962B;
defparam \Add1~56 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N26
cycloneive_lcell_comb \Add1~58 (
// Equation(s):
// \Add1~58_combout  = (\Mux66~0_combout  & ((\Mux2~1_combout  & (!\Add1~57 )) # (!\Mux2~1_combout  & ((\Add1~57 ) # (GND))))) # (!\Mux66~0_combout  & ((\Mux2~1_combout  & (\Add1~57  & VCC)) # (!\Mux2~1_combout  & (!\Add1~57 ))))
// \Add1~59  = CARRY((\Mux66~0_combout  & ((!\Add1~57 ) # (!\Mux2~1_combout ))) # (!\Mux66~0_combout  & (!\Mux2~1_combout  & !\Add1~57 )))

	.dataa(Mux66),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~57 ),
	.combout(\Add1~58_combout ),
	.cout(\Add1~59 ));
// synopsys translate_off
defparam \Add1~58 .lut_mask = 16'h692B;
defparam \Add1~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N14
cycloneive_lcell_comb \aluif.portOut[29]~164 (
// Equation(s):
// \aluif.portOut[29]~164_combout  = (\aluif.portOut[2]~32_combout  & (\aluif.portOut[5]~25_combout  & (\Mux66~0_combout  $ (\Mux2~1_combout ))))

	.dataa(\aluif.portOut[2]~32_combout ),
	.datab(Mux66),
	.datac(Mux2),
	.datad(\aluif.portOut[5]~25_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[29]~164_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~164 .lut_mask = 16'h2800;
defparam \aluif.portOut[29]~164 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N8
cycloneive_lcell_comb \portOut~52 (
// Equation(s):
// \portOut~52_combout  = (\Mux66~0_combout ) # (\Mux2~1_combout )

	.dataa(gnd),
	.datab(Mux66),
	.datac(gnd),
	.datad(Mux2),
	.cin(gnd),
	.combout(\portOut~52_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~52 .lut_mask = 16'hFFCC;
defparam \portOut~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N6
cycloneive_lcell_comb \aluif.portOut[29]~155 (
// Equation(s):
// \aluif.portOut[29]~155_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & (\ShiftRight0~109_combout )) # (!\prif.ALUOP_ex [2] & ((\portOut~52_combout ))))) # (!\aluif.portOut[15]~26_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\ShiftRight0~109_combout ),
	.datab(\aluif.portOut[15]~26_combout ),
	.datac(\portOut~52_combout ),
	.datad(prifALUOP_ex_2),
	.cin(gnd),
	.combout(\aluif.portOut[29]~155_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~155 .lut_mask = 16'h88F3;
defparam \aluif.portOut[29]~155 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N26
cycloneive_lcell_comb \aluif.portOut[29]~163 (
// Equation(s):
// \aluif.portOut[29]~163_combout  = (!\prif.ALUOP_ex [0] & ((\prif.ALUOP_ex [1] & ((\aluif.portOut[29]~155_combout ))) # (!\prif.ALUOP_ex [1] & ((!\aluif.portOut[29]~155_combout ) # (!\portOut~52_combout )))))

	.dataa(prifALUOP_ex_0),
	.datab(\portOut~52_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.portOut[29]~155_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[29]~163_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~163 .lut_mask = 16'h5105;
defparam \aluif.portOut[29]~163 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N16
cycloneive_lcell_comb \aluif.portOut[29]~165 (
// Equation(s):
// \aluif.portOut[29]~165_combout  = (\aluif.portOut[29]~164_combout ) # ((\Add1~58_combout  & (\prif.ALUOP_ex [3] & \aluif.portOut[29]~163_combout )))

	.dataa(\Add1~58_combout ),
	.datab(\aluif.portOut[29]~164_combout ),
	.datac(prifALUOP_ex_3),
	.datad(\aluif.portOut[29]~163_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[29]~165_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~165 .lut_mask = 16'hECCC;
defparam \aluif.portOut[29]~165 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N22
cycloneive_lcell_comb \ShiftLeft0~88 (
// Equation(s):
// \ShiftLeft0~88_combout  = (\Mux95~1_combout  & (\Mux5~1_combout )) # (!\Mux95~1_combout  & ((\Mux4~1_combout )))

	.dataa(Mux95),
	.datab(Mux5),
	.datac(gnd),
	.datad(Mux4),
	.cin(gnd),
	.combout(\ShiftLeft0~88_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~88 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N28
cycloneive_lcell_comb \aluif.portOut[29]~158 (
// Equation(s):
// \aluif.portOut[29]~158_combout  = (\aluif.portOut[29]~157_combout  & (((\ShiftLeft0~87_combout ) # (!\aluif.portOut[2]~35_combout )))) # (!\aluif.portOut[29]~157_combout  & (\ShiftLeft0~88_combout  & ((\aluif.portOut[2]~35_combout ))))

	.dataa(\aluif.portOut[29]~157_combout ),
	.datab(\ShiftLeft0~88_combout ),
	.datac(\ShiftLeft0~87_combout ),
	.datad(\aluif.portOut[2]~35_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[29]~158_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~158 .lut_mask = 16'hE4AA;
defparam \aluif.portOut[29]~158 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N6
cycloneive_lcell_comb \aluif.portOut[29]~159 (
// Equation(s):
// \aluif.portOut[29]~159_combout  = (\aluif.portOut[1]~13_combout  & ((\aluif.portOut[2]~34_combout  & ((\ShiftLeft0~57_combout ))) # (!\aluif.portOut[2]~34_combout  & (\aluif.portOut[29]~158_combout )))) # (!\aluif.portOut[1]~13_combout  & 
// (((\aluif.portOut[2]~34_combout ))))

	.dataa(\aluif.portOut[1]~13_combout ),
	.datab(\aluif.portOut[29]~158_combout ),
	.datac(\aluif.portOut[2]~34_combout ),
	.datad(\ShiftLeft0~57_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[29]~159_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~159 .lut_mask = 16'hF858;
defparam \aluif.portOut[29]~159 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N16
cycloneive_lcell_comb \Add0~48 (
// Equation(s):
// \Add0~48_combout  = ((\Mux71~0_combout  $ (\Mux7~1_combout  $ (!\Add0~47 )))) # (GND)
// \Add0~49  = CARRY((\Mux71~0_combout  & ((\Mux7~1_combout ) # (!\Add0~47 ))) # (!\Mux71~0_combout  & (\Mux7~1_combout  & !\Add0~47 )))

	.dataa(Mux71),
	.datab(Mux7),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~47 ),
	.combout(\Add0~48_combout ),
	.cout(\Add0~49 ));
// synopsys translate_off
defparam \Add0~48 .lut_mask = 16'h698E;
defparam \Add0~48 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N18
cycloneive_lcell_comb \Add0~50 (
// Equation(s):
// \Add0~50_combout  = (\Mux70~0_combout  & ((\Mux6~1_combout  & (\Add0~49  & VCC)) # (!\Mux6~1_combout  & (!\Add0~49 )))) # (!\Mux70~0_combout  & ((\Mux6~1_combout  & (!\Add0~49 )) # (!\Mux6~1_combout  & ((\Add0~49 ) # (GND)))))
// \Add0~51  = CARRY((\Mux70~0_combout  & (!\Mux6~1_combout  & !\Add0~49 )) # (!\Mux70~0_combout  & ((!\Add0~49 ) # (!\Mux6~1_combout ))))

	.dataa(Mux70),
	.datab(Mux6),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~49 ),
	.combout(\Add0~50_combout ),
	.cout(\Add0~51 ));
// synopsys translate_off
defparam \Add0~50 .lut_mask = 16'h9617;
defparam \Add0~50 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N20
cycloneive_lcell_comb \Add0~52 (
// Equation(s):
// \Add0~52_combout  = ((\Mux5~1_combout  $ (\Mux69~0_combout  $ (!\Add0~51 )))) # (GND)
// \Add0~53  = CARRY((\Mux5~1_combout  & ((\Mux69~0_combout ) # (!\Add0~51 ))) # (!\Mux5~1_combout  & (\Mux69~0_combout  & !\Add0~51 )))

	.dataa(Mux5),
	.datab(Mux69),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~51 ),
	.combout(\Add0~52_combout ),
	.cout(\Add0~53 ));
// synopsys translate_off
defparam \Add0~52 .lut_mask = 16'h698E;
defparam \Add0~52 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N22
cycloneive_lcell_comb \Add0~54 (
// Equation(s):
// \Add0~54_combout  = (\Mux68~0_combout  & ((\Mux4~1_combout  & (\Add0~53  & VCC)) # (!\Mux4~1_combout  & (!\Add0~53 )))) # (!\Mux68~0_combout  & ((\Mux4~1_combout  & (!\Add0~53 )) # (!\Mux4~1_combout  & ((\Add0~53 ) # (GND)))))
// \Add0~55  = CARRY((\Mux68~0_combout  & (!\Mux4~1_combout  & !\Add0~53 )) # (!\Mux68~0_combout  & ((!\Add0~53 ) # (!\Mux4~1_combout ))))

	.dataa(Mux68),
	.datab(Mux4),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~53 ),
	.combout(\Add0~54_combout ),
	.cout(\Add0~55 ));
// synopsys translate_off
defparam \Add0~54 .lut_mask = 16'h9617;
defparam \Add0~54 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N26
cycloneive_lcell_comb \Add0~58 (
// Equation(s):
// \Add0~58_combout  = (\Mux66~0_combout  & ((\Mux2~1_combout  & (\Add0~57  & VCC)) # (!\Mux2~1_combout  & (!\Add0~57 )))) # (!\Mux66~0_combout  & ((\Mux2~1_combout  & (!\Add0~57 )) # (!\Mux2~1_combout  & ((\Add0~57 ) # (GND)))))
// \Add0~59  = CARRY((\Mux66~0_combout  & (!\Mux2~1_combout  & !\Add0~57 )) # (!\Mux66~0_combout  & ((!\Add0~57 ) # (!\Mux2~1_combout ))))

	.dataa(Mux66),
	.datab(Mux2),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~57 ),
	.combout(\Add0~58_combout ),
	.cout(\Add0~59 ));
// synopsys translate_off
defparam \Add0~58 .lut_mask = 16'h9617;
defparam \Add0~58 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N0
cycloneive_lcell_comb \aluif.portOut[29]~160 (
// Equation(s):
// \aluif.portOut[29]~160_combout  = (\aluif.portOut[1]~13_combout  & (((\aluif.portOut[29]~159_combout )))) # (!\aluif.portOut[1]~13_combout  & (\Mux2~1_combout  & (\Mux66~0_combout  & !\aluif.portOut[29]~159_combout )))

	.dataa(\aluif.portOut[1]~13_combout ),
	.datab(Mux2),
	.datac(Mux66),
	.datad(\aluif.portOut[29]~159_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[29]~160_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~160 .lut_mask = 16'hAA40;
defparam \aluif.portOut[29]~160 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N4
cycloneive_lcell_comb \aluif.portOut[29]~162 (
// Equation(s):
// \aluif.portOut[29]~162_combout  = (\Add0~58_combout  & ((\aluif.portOut[29]~159_combout ) # ((\aluif.portOut[29]~160_combout )))) # (!\Add0~58_combout  & (((\Add1~58_combout  & \aluif.portOut[29]~160_combout ))))

	.dataa(\aluif.portOut[29]~159_combout ),
	.datab(\Add0~58_combout ),
	.datac(\Add1~58_combout ),
	.datad(\aluif.portOut[29]~160_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[29]~162_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~162 .lut_mask = 16'hFC88;
defparam \aluif.portOut[29]~162 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y24_N28
cycloneive_lcell_comb \aluif.portOut[29]~156 (
// Equation(s):
// \aluif.portOut[29]~156_combout  = (!\prif.ALUOP_ex [0] & (\prif.ALUOP_ex [3] & ((\prif.ALUOP_ex [1]) # (!\portOut~52_combout ))))

	.dataa(prifALUOP_ex_0),
	.datab(prifALUOP_ex_1),
	.datac(\portOut~52_combout ),
	.datad(prifALUOP_ex_3),
	.cin(gnd),
	.combout(\aluif.portOut[29]~156_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~156 .lut_mask = 16'h4500;
defparam \aluif.portOut[29]~156 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y23_N10
cycloneive_lcell_comb \aluif.portOut[29]~161 (
// Equation(s):
// \aluif.portOut[29]~161_combout  = (\aluif.portOut[29]~155_combout  & ((\aluif.portOut[29]~156_combout ) # ((\aluif.portOut[28]~154_combout  & \aluif.portOut[29]~160_combout )))) # (!\aluif.portOut[29]~155_combout  & (((\aluif.portOut[28]~154_combout  & 
// \aluif.portOut[29]~160_combout ))))

	.dataa(\aluif.portOut[29]~155_combout ),
	.datab(\aluif.portOut[29]~156_combout ),
	.datac(\aluif.portOut[28]~154_combout ),
	.datad(\aluif.portOut[29]~160_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[29]~161_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[29]~161 .lut_mask = 16'hF888;
defparam \aluif.portOut[29]~161 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N2
cycloneive_lcell_comb \aluif.portOut[28]~168 (
// Equation(s):
// \aluif.portOut[28]~168_combout  = (\Mux3~1_combout ) # (\Mux67~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux3),
	.datad(Mux67),
	.cin(gnd),
	.combout(\aluif.portOut[28]~168_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~168 .lut_mask = 16'hFFF0;
defparam \aluif.portOut[28]~168 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N4
cycloneive_lcell_comb \aluif.portOut[28]~171 (
// Equation(s):
// \aluif.portOut[28]~171_combout  = (\prif.ALUOP_ex [2] & (((\ShiftRight0~110_combout  & \aluif.portOut[15]~26_combout )))) # (!\prif.ALUOP_ex [2] & ((\aluif.portOut[28]~168_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\aluif.portOut[28]~168_combout ),
	.datac(\ShiftRight0~110_combout ),
	.datad(\aluif.portOut[15]~26_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~171_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~171 .lut_mask = 16'hE455;
defparam \aluif.portOut[28]~171 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N10
cycloneive_lcell_comb \aluif.portOut[28]~262 (
// Equation(s):
// \aluif.portOut[28]~262_combout  = (\aluif.portOut[28]~171_combout  & ((\prif.ALUOP_ex [1]) # ((!\Mux67~0_combout  & !\Mux3~1_combout ))))

	.dataa(Mux67),
	.datab(Mux3),
	.datac(\aluif.portOut[28]~171_combout ),
	.datad(prifALUOP_ex_1),
	.cin(gnd),
	.combout(\aluif.portOut[28]~262_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~262 .lut_mask = 16'hF010;
defparam \aluif.portOut[28]~262 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N6
cycloneive_lcell_comb \ShiftLeft0~92 (
// Equation(s):
// \ShiftLeft0~92_combout  = (\Mux95~1_combout  & ((\Mux6~1_combout ))) # (!\Mux95~1_combout  & (\Mux5~1_combout ))

	.dataa(gnd),
	.datab(Mux5),
	.datac(Mux95),
	.datad(Mux6),
	.cin(gnd),
	.combout(\ShiftLeft0~92_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~92 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N6
cycloneive_lcell_comb \ShiftLeft0~96 (
// Equation(s):
// \ShiftLeft0~96_combout  = (\Mux94~1_combout  & (((\Mux95~1_combout ) # (\Mux13~1_combout )))) # (!\Mux94~1_combout  & (\Mux11~1_combout  & (!\Mux95~1_combout )))

	.dataa(Mux11),
	.datab(Mux94),
	.datac(Mux95),
	.datad(Mux13),
	.cin(gnd),
	.combout(\ShiftLeft0~96_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~96 .lut_mask = 16'hCEC2;
defparam \ShiftLeft0~96 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N8
cycloneive_lcell_comb \ShiftLeft0~97 (
// Equation(s):
// \ShiftLeft0~97_combout  = (\Mux95~1_combout  & ((\ShiftLeft0~96_combout  & ((\Mux14~1_combout ))) # (!\ShiftLeft0~96_combout  & (\Mux12~1_combout )))) # (!\Mux95~1_combout  & (((\ShiftLeft0~96_combout ))))

	.dataa(Mux95),
	.datab(Mux12),
	.datac(Mux14),
	.datad(\ShiftLeft0~96_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~97_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~97 .lut_mask = 16'hF588;
defparam \ShiftLeft0~97 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y22_N14
cycloneive_lcell_comb \ShiftLeft0~99 (
// Equation(s):
// \ShiftLeft0~99_combout  = (!\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux16~1_combout ))) # (!\Mux95~1_combout  & (\Mux15~1_combout ))))

	.dataa(Mux94),
	.datab(Mux95),
	.datac(Mux15),
	.datad(Mux16),
	.cin(gnd),
	.combout(\ShiftLeft0~99_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~99 .lut_mask = 16'h5410;
defparam \ShiftLeft0~99 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N26
cycloneive_lcell_comb \ShiftLeft0~100 (
// Equation(s):
// \ShiftLeft0~100_combout  = (\Mux93~2_combout  & ((\ShiftLeft0~98_combout ) # ((\ShiftLeft0~99_combout )))) # (!\Mux93~2_combout  & (((\ShiftLeft0~97_combout ))))

	.dataa(\ShiftLeft0~98_combout ),
	.datab(Mux931),
	.datac(\ShiftLeft0~97_combout ),
	.datad(\ShiftLeft0~99_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~100_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~100 .lut_mask = 16'hFCB8;
defparam \ShiftLeft0~100 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N24
cycloneive_lcell_comb \aluif.portOut[28]~174 (
// Equation(s):
// \aluif.portOut[28]~174_combout  = (\aluif.portOut[28]~173_combout  & (((\ShiftLeft0~100_combout ) # (!\aluif.portOut[2]~35_combout )))) # (!\aluif.portOut[28]~173_combout  & (\ShiftLeft0~92_combout  & (\aluif.portOut[2]~35_combout )))

	.dataa(\aluif.portOut[28]~173_combout ),
	.datab(\ShiftLeft0~92_combout ),
	.datac(\aluif.portOut[2]~35_combout ),
	.datad(\ShiftLeft0~100_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~174_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~174 .lut_mask = 16'hEA4A;
defparam \aluif.portOut[28]~174 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N18
cycloneive_lcell_comb \aluif.portOut[28]~177 (
// Equation(s):
// \aluif.portOut[28]~177_combout  = (\aluif.portOut[1]~13_combout  & (((\aluif.portOut[28]~174_combout ) # (\aluif.portOut[2]~34_combout )))) # (!\aluif.portOut[1]~13_combout  & (\portOut~53_combout  & ((!\aluif.portOut[2]~34_combout ))))

	.dataa(\portOut~53_combout ),
	.datab(\aluif.portOut[1]~13_combout ),
	.datac(\aluif.portOut[28]~174_combout ),
	.datad(\aluif.portOut[2]~34_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~177_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~177 .lut_mask = 16'hCCE2;
defparam \aluif.portOut[28]~177 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N26
cycloneive_lcell_comb \portOut~53 (
// Equation(s):
// \portOut~53_combout  = (\Mux3~1_combout  & \Mux67~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux3),
	.datad(Mux67),
	.cin(gnd),
	.combout(\portOut~53_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~53 .lut_mask = 16'hF000;
defparam \portOut~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N0
cycloneive_lcell_comb \aluif.portOut[28]~172 (
// Equation(s):
// \aluif.portOut[28]~172_combout  = (\aluif.portOut[28]~170_combout  & (\aluif.portOut[28]~171_combout  & ((\prif.ALUOP_ex [1]) # (!\aluif.portOut[28]~168_combout ))))

	.dataa(\aluif.portOut[28]~170_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\aluif.portOut[28]~171_combout ),
	.datad(\aluif.portOut[28]~168_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~172_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~172 .lut_mask = 16'h80A0;
defparam \aluif.portOut[28]~172 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N24
cycloneive_lcell_comb \aluif.portOut[28]~176 (
// Equation(s):
// \aluif.portOut[28]~176_combout  = (\aluif.portOut[28]~175_combout ) # ((\aluif.portOut[28]~172_combout ) # ((!\aluif.portOut[1]~13_combout  & \portOut~53_combout )))

	.dataa(\aluif.portOut[28]~175_combout ),
	.datab(\aluif.portOut[1]~13_combout ),
	.datac(\portOut~53_combout ),
	.datad(\aluif.portOut[28]~172_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~176_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~176 .lut_mask = 16'hFFBA;
defparam \aluif.portOut[28]~176 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N16
cycloneive_lcell_comb \aluif.portOut[28]~178 (
// Equation(s):
// \aluif.portOut[28]~178_combout  = (\aluif.portOut[28]~154_combout  & ((\Add0~56_combout ) # ((\aluif.portOut[28]~177_combout ) # (!\aluif.portOut[28]~176_combout ))))

	.dataa(\Add0~56_combout ),
	.datab(\aluif.portOut[28]~177_combout ),
	.datac(\aluif.portOut[28]~154_combout ),
	.datad(\aluif.portOut[28]~176_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~178_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~178 .lut_mask = 16'hE0F0;
defparam \aluif.portOut[28]~178 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N8
cycloneive_lcell_comb \aluif.portOut[28]~169 (
// Equation(s):
// \aluif.portOut[28]~169_combout  = (\prif.ALUOP_ex [2] & (((\ShiftRight0~110_combout  & \aluif.portOut[15]~26_combout )))) # (!\prif.ALUOP_ex [2] & ((\aluif.portOut[28]~168_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\aluif.portOut[28]~168_combout ),
	.datac(\ShiftRight0~110_combout ),
	.datad(\aluif.portOut[15]~26_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~169_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~169 .lut_mask = 16'hE455;
defparam \aluif.portOut[28]~169 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N30
cycloneive_lcell_comb \aluif.portOut[28]~170 (
// Equation(s):
// \aluif.portOut[28]~170_combout  = (aluifportOut_5 & ((\prif.ALUOP_ex [1] & (\aluif.portOut[28]~169_combout )) # (!\prif.ALUOP_ex [1] & ((!\aluif.portOut[28]~168_combout ) # (!\aluif.portOut[28]~169_combout )))))

	.dataa(aluifportOut_5),
	.datab(prifALUOP_ex_1),
	.datac(\aluif.portOut[28]~169_combout ),
	.datad(\aluif.portOut[28]~168_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~170_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~170 .lut_mask = 16'h82A2;
defparam \aluif.portOut[28]~170 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N22
cycloneive_lcell_comb \aluif.portOut[28]~179 (
// Equation(s):
// \aluif.portOut[28]~179_combout  = (\aluif.portOut[28]~178_combout  & (((\aluif.portOut[28]~176_combout )))) # (!\aluif.portOut[28]~178_combout  & (\aluif.portOut[28]~262_combout  & (\aluif.portOut[28]~170_combout )))

	.dataa(\aluif.portOut[28]~262_combout ),
	.datab(\aluif.portOut[28]~178_combout ),
	.datac(\aluif.portOut[28]~170_combout ),
	.datad(\aluif.portOut[28]~176_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[28]~179_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~179 .lut_mask = 16'hEC20;
defparam \aluif.portOut[28]~179 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y21_N20
cycloneive_lcell_comb \aluif.portOut[28]~167 (
// Equation(s):
// \aluif.portOut[28]~167_combout  = (\aluif.portOut[2]~32_combout  & (\aluif.portOut[5]~25_combout  & (\Mux3~1_combout  $ (\Mux67~0_combout ))))

	.dataa(\aluif.portOut[2]~32_combout ),
	.datab(\aluif.portOut[5]~25_combout ),
	.datac(Mux3),
	.datad(Mux67),
	.cin(gnd),
	.combout(\aluif.portOut[28]~167_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[28]~167 .lut_mask = 16'h0880;
defparam \aluif.portOut[28]~167 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N28
cycloneive_lcell_comb \Add0~60 (
// Equation(s):
// \Add0~60_combout  = ((\Mux1~1_combout  $ (\Mux65~0_combout  $ (!\Add0~59 )))) # (GND)
// \Add0~61  = CARRY((\Mux1~1_combout  & ((\Mux65~0_combout ) # (!\Add0~59 ))) # (!\Mux1~1_combout  & (\Mux65~0_combout  & !\Add0~59 )))

	.dataa(Mux1),
	.datab(Mux65),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add0~59 ),
	.combout(\Add0~60_combout ),
	.cout(\Add0~61 ));
// synopsys translate_off
defparam \Add0~60 .lut_mask = 16'h698E;
defparam \Add0~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X55_Y24_N30
cycloneive_lcell_comb \Add0~62 (
// Equation(s):
// \Add0~62_combout  = \Mux0~1_combout  $ (\Add0~61  $ (\Mux64~0_combout ))

	.dataa(gnd),
	.datab(Mux0),
	.datac(gnd),
	.datad(Mux64),
	.cin(\Add0~61 ),
	.combout(\Add0~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~62 .lut_mask = 16'hC33C;
defparam \Add0~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N28
cycloneive_lcell_comb \Add1~60 (
// Equation(s):
// \Add1~60_combout  = ((\Mux65~0_combout  $ (\Mux1~1_combout  $ (\Add1~59 )))) # (GND)
// \Add1~61  = CARRY((\Mux65~0_combout  & (\Mux1~1_combout  & !\Add1~59 )) # (!\Mux65~0_combout  & ((\Mux1~1_combout ) # (!\Add1~59 ))))

	.dataa(Mux65),
	.datab(Mux1),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~59 ),
	.combout(\Add1~60_combout ),
	.cout(\Add1~61 ));
// synopsys translate_off
defparam \Add1~60 .lut_mask = 16'h964D;
defparam \Add1~60 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X58_Y24_N30
cycloneive_lcell_comb \Add1~62 (
// Equation(s):
// \Add1~62_combout  = \Mux0~1_combout  $ (\Add1~61  $ (!\Mux64~0_combout ))

	.dataa(gnd),
	.datab(Mux0),
	.datac(gnd),
	.datad(Mux64),
	.cin(\Add1~61 ),
	.combout(\Add1~62_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~62 .lut_mask = 16'h3CC3;
defparam \Add1~62 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N2
cycloneive_lcell_comb \portOut~54 (
// Equation(s):
// \portOut~54_combout  = (\Mux64~0_combout ) # (\Mux0~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux64),
	.datad(Mux0),
	.cin(gnd),
	.combout(\portOut~54_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~54 .lut_mask = 16'hFFF0;
defparam \portOut~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N20
cycloneive_lcell_comb \aluif.neg_flag~12 (
// Equation(s):
// \aluif.neg_flag~12_combout  = (\prif.ALUOP_ex [2] & (\ShiftRight0~113_combout  & (\aluif.portOut[15]~26_combout ))) # (!\prif.ALUOP_ex [2] & (((\portOut~54_combout ) # (!\aluif.portOut[15]~26_combout ))))

	.dataa(\ShiftRight0~113_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\portOut~54_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~12_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~12 .lut_mask = 16'hB383;
defparam \aluif.neg_flag~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N22
cycloneive_lcell_comb \aluif.neg_flag~21 (
// Equation(s):
// \aluif.neg_flag~21_combout  = (\prif.ALUOP_ex [1] & (((\aluif.neg_flag~12_combout )))) # (!\prif.ALUOP_ex [1] & (((!\Mux0~1_combout  & !\Mux64~0_combout )) # (!\aluif.neg_flag~12_combout )))

	.dataa(Mux0),
	.datab(prifALUOP_ex_1),
	.datac(Mux64),
	.datad(\aluif.neg_flag~12_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~21_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~21 .lut_mask = 16'hCD33;
defparam \aluif.neg_flag~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N0
cycloneive_lcell_comb \ShiftLeft0~101 (
// Equation(s):
// \ShiftLeft0~101_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux7~1_combout ))) # (!\Mux95~1_combout  & (\Mux6~1_combout ))))

	.dataa(Mux95),
	.datab(Mux94),
	.datac(Mux6),
	.datad(Mux7),
	.cin(gnd),
	.combout(\ShiftLeft0~101_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~101 .lut_mask = 16'hC840;
defparam \ShiftLeft0~101 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N10
cycloneive_lcell_comb \ShiftLeft0~102 (
// Equation(s):
// \ShiftLeft0~102_combout  = (\ShiftLeft0~101_combout ) # ((\ShiftLeft0~88_combout  & !\Mux94~1_combout ))

	.dataa(\ShiftLeft0~88_combout ),
	.datab(gnd),
	.datac(Mux94),
	.datad(\ShiftLeft0~101_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~102_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~102 .lut_mask = 16'hFF0A;
defparam \ShiftLeft0~102 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N22
cycloneive_lcell_comb \aluif.portOut[30]~181 (
// Equation(s):
// \aluif.portOut[30]~181_combout  = (\Mux93~2_combout ) # ((\Mux95~1_combout  & !\Mux94~1_combout ))

	.dataa(Mux931),
	.datab(gnd),
	.datac(Mux95),
	.datad(Mux94),
	.cin(gnd),
	.combout(\aluif.portOut[30]~181_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[30]~181 .lut_mask = 16'hAAFA;
defparam \aluif.portOut[30]~181 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N0
cycloneive_lcell_comb \ShiftLeft0~91 (
// Equation(s):
// \ShiftLeft0~91_combout  = (\Mux95~1_combout  & ((\Mux3~1_combout ))) # (!\Mux95~1_combout  & (\Mux2~1_combout ))

	.dataa(gnd),
	.datab(Mux2),
	.datac(Mux3),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftLeft0~91_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~91 .lut_mask = 16'hF0CC;
defparam \ShiftLeft0~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N12
cycloneive_lcell_comb \aluif.neg_flag~14 (
// Equation(s):
// \aluif.neg_flag~14_combout  = (\ShiftLeft0~5_combout  & (((\aluif.portOut[30]~181_combout ) # (\ShiftLeft0~91_combout )))) # (!\ShiftLeft0~5_combout  & (\Mux0~1_combout  & (!\aluif.portOut[30]~181_combout )))

	.dataa(Mux0),
	.datab(\ShiftLeft0~5_combout ),
	.datac(\aluif.portOut[30]~181_combout ),
	.datad(\ShiftLeft0~91_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~14_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~14 .lut_mask = 16'hCEC2;
defparam \aluif.neg_flag~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y23_N14
cycloneive_lcell_comb \aluif.neg_flag~15 (
// Equation(s):
// \aluif.neg_flag~15_combout  = (\aluif.portOut[30]~181_combout  & ((\aluif.neg_flag~14_combout  & ((\ShiftLeft0~102_combout ))) # (!\aluif.neg_flag~14_combout  & (\Mux1~1_combout )))) # (!\aluif.portOut[30]~181_combout  & (((\aluif.neg_flag~14_combout ))))

	.dataa(\aluif.portOut[30]~181_combout ),
	.datab(Mux1),
	.datac(\ShiftLeft0~102_combout ),
	.datad(\aluif.neg_flag~14_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~15_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~15 .lut_mask = 16'hF588;
defparam \aluif.neg_flag~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N24
cycloneive_lcell_comb \aluif.neg_flag~16 (
// Equation(s):
// \aluif.neg_flag~16_combout  = (\aluif.neg_flag~13_combout  & (((\ShiftLeft0~77_combout ) # (\aluif.portOut[15]~81_combout )))) # (!\aluif.neg_flag~13_combout  & (\aluif.neg_flag~15_combout  & ((!\aluif.portOut[15]~81_combout ))))

	.dataa(\aluif.neg_flag~13_combout ),
	.datab(\aluif.neg_flag~15_combout ),
	.datac(\ShiftLeft0~77_combout ),
	.datad(\aluif.portOut[15]~81_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~16_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~16 .lut_mask = 16'hAAE4;
defparam \aluif.neg_flag~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N16
cycloneive_lcell_comb \aluif.neg_flag~18 (
// Equation(s):
// \aluif.neg_flag~18_combout  = (\aluif.portOut[23]~135_combout  & (!\aluif.portOut[23]~136_combout  & (\aluif.neg_flag~21_combout ))) # (!\aluif.portOut[23]~135_combout  & ((\aluif.portOut[23]~136_combout ) # ((\aluif.neg_flag~16_combout ))))

	.dataa(\aluif.portOut[23]~135_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(\aluif.neg_flag~21_combout ),
	.datad(\aluif.neg_flag~16_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~18_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~18 .lut_mask = 16'h7564;
defparam \aluif.neg_flag~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N8
cycloneive_lcell_comb \aluif.neg_flag~20 (
// Equation(s):
// \aluif.neg_flag~20_combout  = (\aluif.neg_flag~12_combout  & ((\prif.ALUOP_ex [1]) # ((!\Mux0~1_combout  & !\Mux64~0_combout ))))

	.dataa(Mux0),
	.datab(prifALUOP_ex_1),
	.datac(Mux64),
	.datad(\aluif.neg_flag~12_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~20_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~20 .lut_mask = 16'hCD00;
defparam \aluif.neg_flag~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N6
cycloneive_lcell_comb \aluif.neg_flag~17 (
// Equation(s):
// \aluif.neg_flag~17_combout  = (\aluif.neg_flag~23_combout  & (!\aluif.portOut[23]~136_combout  & (\aluif.neg_flag~20_combout ))) # (!\aluif.neg_flag~23_combout  & ((\aluif.portOut[23]~136_combout ) # ((\aluif.neg_flag~16_combout ))))

	.dataa(\aluif.neg_flag~23_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(\aluif.neg_flag~20_combout ),
	.datad(\aluif.neg_flag~16_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~17_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~17 .lut_mask = 16'h7564;
defparam \aluif.neg_flag~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N4
cycloneive_lcell_comb \aluif.neg_flag~22 (
// Equation(s):
// \aluif.neg_flag~22_combout  = (\prif.ALUOP_ex [0] & ((\aluif.neg_flag~18_combout  & (\prif.ALUOP_ex [1])) # (!\aluif.neg_flag~18_combout  & (!\prif.ALUOP_ex [1] & \aluif.neg_flag~17_combout )))) # (!\prif.ALUOP_ex [0] & (\aluif.neg_flag~18_combout ))

	.dataa(prifALUOP_ex_0),
	.datab(\aluif.neg_flag~18_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.neg_flag~17_combout ),
	.cin(gnd),
	.combout(\aluif.neg_flag~22_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.neg_flag~22 .lut_mask = 16'hC6C4;
defparam \aluif.neg_flag~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N18
cycloneive_lcell_comb \portOut~59 (
// Equation(s):
// \portOut~59_combout  = \Mux65~0_combout  $ (\Mux1~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux65),
	.datad(Mux1),
	.cin(gnd),
	.combout(\portOut~59_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~59 .lut_mask = 16'h0FF0;
defparam \portOut~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N28
cycloneive_lcell_comb \portOut~57 (
// Equation(s):
// \portOut~57_combout  = (\Mux65~0_combout ) # (\Mux1~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux65),
	.datad(Mux1),
	.cin(gnd),
	.combout(\portOut~57_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~57 .lut_mask = 16'hFFF0;
defparam \portOut~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N26
cycloneive_lcell_comb \aluif.portOut[30]~182 (
// Equation(s):
// \aluif.portOut[30]~182_combout  = (\prif.ALUOP_ex [2] & (\ShiftRight0~111_combout  & (\aluif.portOut[15]~26_combout ))) # (!\prif.ALUOP_ex [2] & (((\portOut~57_combout ) # (!\aluif.portOut[15]~26_combout ))))

	.dataa(\ShiftRight0~111_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\portOut~57_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[30]~182_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[30]~182 .lut_mask = 16'hB383;
defparam \aluif.portOut[30]~182 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N0
cycloneive_lcell_comb \aluif.portOut[30]~183 (
// Equation(s):
// \aluif.portOut[30]~183_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[30]~182_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[30]~182_combout  & ((!\portOut~57_combout ))) # (!\aluif.portOut[30]~182_combout  & (\Add1~60_combout ))))

	.dataa(\Add1~60_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\aluif.portOut[30]~182_combout ),
	.datad(\portOut~57_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[30]~183_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[30]~183 .lut_mask = 16'hC2F2;
defparam \aluif.portOut[30]~183 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N26
cycloneive_lcell_comb \ShiftLeft0~68 (
// Equation(s):
// \ShiftLeft0~68_combout  = (\Mux92~2_combout  & ((\Mux93~2_combout  & (\ShiftLeft0~21_combout )) # (!\Mux93~2_combout  & ((\ShiftLeft0~35_combout )))))

	.dataa(Mux92),
	.datab(\ShiftLeft0~21_combout ),
	.datac(Mux931),
	.datad(\ShiftLeft0~35_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~68_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~68 .lut_mask = 16'h8A80;
defparam \ShiftLeft0~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N14
cycloneive_lcell_comb \ShiftLeft0~72 (
// Equation(s):
// \ShiftLeft0~72_combout  = (\ShiftLeft0~68_combout ) # ((!\Mux92~2_combout  & \ShiftLeft0~71_combout ))

	.dataa(Mux92),
	.datab(gnd),
	.datac(\ShiftLeft0~68_combout ),
	.datad(\ShiftLeft0~71_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~72_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~72 .lut_mask = 16'hF5F0;
defparam \ShiftLeft0~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y22_N24
cycloneive_lcell_comb \aluif.portOut[30]~186 (
// Equation(s):
// \aluif.portOut[30]~186_combout  = (\aluif.portOut[15]~82_combout  & ((\aluif.portOut[15]~83_combout  & (\portOut~58_combout )) # (!\aluif.portOut[15]~83_combout  & ((\ShiftLeft0~72_combout ))))) # (!\aluif.portOut[15]~82_combout  & 
// (((\aluif.portOut[15]~83_combout ))))

	.dataa(\portOut~58_combout ),
	.datab(\aluif.portOut[15]~82_combout ),
	.datac(\aluif.portOut[15]~83_combout ),
	.datad(\ShiftLeft0~72_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[30]~186_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[30]~186 .lut_mask = 16'hBCB0;
defparam \aluif.portOut[30]~186 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N24
cycloneive_lcell_comb \aluif.portOut[30]~187 (
// Equation(s):
// \aluif.portOut[30]~187_combout  = (\aluif.portOut[30]~186_combout  & (((\ShiftLeft0~82_combout ) # (\aluif.portOut[15]~81_combout )))) # (!\aluif.portOut[30]~186_combout  & (\aluif.portOut[30]~185_combout  & ((!\aluif.portOut[15]~81_combout ))))

	.dataa(\aluif.portOut[30]~185_combout ),
	.datab(\aluif.portOut[30]~186_combout ),
	.datac(\ShiftLeft0~82_combout ),
	.datad(\aluif.portOut[15]~81_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[30]~187_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[30]~187 .lut_mask = 16'hCCE2;
defparam \aluif.portOut[30]~187 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y22_N10
cycloneive_lcell_comb \aluif.portOut[30]~188 (
// Equation(s):
// \aluif.portOut[30]~188_combout  = (\aluif.portOut[23]~135_combout  & (\aluif.portOut[23]~136_combout )) # (!\aluif.portOut[23]~135_combout  & ((\aluif.portOut[23]~136_combout  & (\Add0~60_combout )) # (!\aluif.portOut[23]~136_combout  & 
// ((\aluif.portOut[30]~187_combout )))))

	.dataa(\aluif.portOut[23]~135_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(\Add0~60_combout ),
	.datad(\aluif.portOut[30]~187_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[30]~188_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[30]~188 .lut_mask = 16'hD9C8;
defparam \aluif.portOut[30]~188 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N24
cycloneive_lcell_comb \portOut~62 (
// Equation(s):
// \portOut~62_combout  = \Mux75~0_combout  $ (\Mux11~1_combout )

	.dataa(Mux75),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux11),
	.cin(gnd),
	.combout(\portOut~62_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~62 .lut_mask = 16'h55AA;
defparam \portOut~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N14
cycloneive_lcell_comb \portOut~60 (
// Equation(s):
// \portOut~60_combout  = (\Mux75~0_combout  & \Mux11~1_combout )

	.dataa(Mux75),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux11),
	.cin(gnd),
	.combout(\portOut~60_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~60 .lut_mask = 16'hAA00;
defparam \portOut~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N4
cycloneive_lcell_comb \aluif.portOut[20]~190 (
// Equation(s):
// \aluif.portOut[20]~190_combout  = (\aluif.portOut[15]~82_combout  & ((\aluif.portOut[15]~83_combout  & ((\portOut~60_combout ))) # (!\aluif.portOut[15]~83_combout  & (\ShiftLeft0~29_combout )))) # (!\aluif.portOut[15]~82_combout  & 
// (((\aluif.portOut[15]~83_combout ))))

	.dataa(\ShiftLeft0~29_combout ),
	.datab(\aluif.portOut[15]~82_combout ),
	.datac(\portOut~60_combout ),
	.datad(\aluif.portOut[15]~83_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[20]~190_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[20]~190 .lut_mask = 16'hF388;
defparam \aluif.portOut[20]~190 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N26
cycloneive_lcell_comb \aluif.portOut[20]~191 (
// Equation(s):
// \aluif.portOut[20]~191_combout  = (\aluif.portOut[20]~190_combout  & ((\ShiftLeft0~61_combout ) # ((\aluif.portOut[15]~81_combout )))) # (!\aluif.portOut[20]~190_combout  & (((\ShiftLeft0~100_combout  & !\aluif.portOut[15]~81_combout ))))

	.dataa(\ShiftLeft0~61_combout ),
	.datab(\ShiftLeft0~100_combout ),
	.datac(\aluif.portOut[20]~190_combout ),
	.datad(\aluif.portOut[15]~81_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[20]~191_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[20]~191 .lut_mask = 16'hF0AC;
defparam \aluif.portOut[20]~191 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N16
cycloneive_lcell_comb \portOut~61 (
// Equation(s):
// \portOut~61_combout  = (\Mux75~0_combout ) # (\Mux11~1_combout )

	.dataa(Mux75),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux11),
	.cin(gnd),
	.combout(\portOut~61_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~61 .lut_mask = 16'hFFAA;
defparam \portOut~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N0
cycloneive_lcell_comb \aluif.portOut[20]~193 (
// Equation(s):
// \aluif.portOut[20]~193_combout  = (\aluif.portOut[20]~192_combout  & ((\prif.ALUOP_ex [1]) # ((!\portOut~61_combout )))) # (!\aluif.portOut[20]~192_combout  & (!\prif.ALUOP_ex [1] & (\Add1~40_combout )))

	.dataa(\aluif.portOut[20]~192_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\Add1~40_combout ),
	.datad(\portOut~61_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[20]~193_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[20]~193 .lut_mask = 16'h98BA;
defparam \aluif.portOut[20]~193 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y24_N2
cycloneive_lcell_comb \aluif.portOut[20]~194 (
// Equation(s):
// \aluif.portOut[20]~194_combout  = (\aluif.portOut[23]~136_combout  & (\aluif.portOut[23]~135_combout )) # (!\aluif.portOut[23]~136_combout  & ((\aluif.portOut[23]~135_combout  & ((\aluif.portOut[20]~193_combout ))) # (!\aluif.portOut[23]~135_combout  & 
// (\aluif.portOut[20]~191_combout ))))

	.dataa(\aluif.portOut[23]~136_combout ),
	.datab(\aluif.portOut[23]~135_combout ),
	.datac(\aluif.portOut[20]~191_combout ),
	.datad(\aluif.portOut[20]~193_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[20]~194_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[20]~194 .lut_mask = 16'hDC98;
defparam \aluif.portOut[20]~194 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N4
cycloneive_lcell_comb \portOut~65 (
// Equation(s):
// \portOut~65_combout  = \Mux14~1_combout  $ (\Mux78~0_combout )

	.dataa(Mux14),
	.datab(gnd),
	.datac(Mux78),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~65_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~65 .lut_mask = 16'h5A5A;
defparam \portOut~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y21_N28
cycloneive_lcell_comb \portOut~63 (
// Equation(s):
// \portOut~63_combout  = (\Mux14~1_combout ) # (\Mux78~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux14),
	.datad(Mux78),
	.cin(gnd),
	.combout(\portOut~63_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~63 .lut_mask = 16'hFFF0;
defparam \portOut~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y21_N14
cycloneive_lcell_comb \aluif.portOut[17]~196 (
// Equation(s):
// \aluif.portOut[17]~196_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[15]~26_combout  & \ShiftRight0~31_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~63_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\portOut~63_combout ),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\ShiftRight0~31_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[17]~196_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[17]~196 .lut_mask = 16'hE545;
defparam \aluif.portOut[17]~196 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y21_N8
cycloneive_lcell_comb \aluif.portOut[17]~197 (
// Equation(s):
// \aluif.portOut[17]~197_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[17]~196_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[17]~196_combout  & (!\portOut~63_combout )) # (!\aluif.portOut[17]~196_combout  & ((\Add1~34_combout )))))

	.dataa(prifALUOP_ex_1),
	.datab(\portOut~63_combout ),
	.datac(\aluif.portOut[17]~196_combout ),
	.datad(\Add1~34_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[17]~197_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[17]~197 .lut_mask = 16'hB5B0;
defparam \aluif.portOut[17]~197 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N20
cycloneive_lcell_comb \portOut~64 (
// Equation(s):
// \portOut~64_combout  = (\Mux14~1_combout  & \Mux78~0_combout )

	.dataa(Mux14),
	.datab(gnd),
	.datac(Mux78),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~64_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~64 .lut_mask = 16'hA0A0;
defparam \portOut~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N30
cycloneive_lcell_comb \aluif.portOut[17]~198 (
// Equation(s):
// \aluif.portOut[17]~198_combout  = (\aluif.portOut[15]~83_combout  & ((\portOut~64_combout ) # ((!\aluif.portOut[15]~82_combout )))) # (!\aluif.portOut[15]~83_combout  & (((\ShiftLeft0~6_combout  & \aluif.portOut[15]~82_combout ))))

	.dataa(\aluif.portOut[15]~83_combout ),
	.datab(\portOut~64_combout ),
	.datac(\ShiftLeft0~6_combout ),
	.datad(\aluif.portOut[15]~82_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[17]~198_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[17]~198 .lut_mask = 16'hD8AA;
defparam \aluif.portOut[17]~198 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N22
cycloneive_lcell_comb \ShiftLeft0~105 (
// Equation(s):
// \ShiftLeft0~105_combout  = (\Mux93~2_combout  & (\ShiftLeft0~55_combout )) # (!\Mux93~2_combout  & ((\ShiftLeft0~84_combout )))

	.dataa(gnd),
	.datab(Mux931),
	.datac(\ShiftLeft0~55_combout ),
	.datad(\ShiftLeft0~84_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~105 .lut_mask = 16'hF3C0;
defparam \ShiftLeft0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N0
cycloneive_lcell_comb \aluif.portOut[17]~199 (
// Equation(s):
// \aluif.portOut[17]~199_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[17]~198_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[17]~198_combout  & (\ShiftLeft0~39_combout )) # (!\aluif.portOut[17]~198_combout  & 
// ((\ShiftLeft0~105_combout )))))

	.dataa(\ShiftLeft0~39_combout ),
	.datab(\aluif.portOut[15]~81_combout ),
	.datac(\aluif.portOut[17]~198_combout ),
	.datad(\ShiftLeft0~105_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[17]~199_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[17]~199 .lut_mask = 16'hE3E0;
defparam \aluif.portOut[17]~199 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N2
cycloneive_lcell_comb \aluif.portOut[17]~200 (
// Equation(s):
// \aluif.portOut[17]~200_combout  = (\aluif.portOut[23]~135_combout  & ((\aluif.portOut[23]~136_combout ) # ((\aluif.portOut[17]~197_combout )))) # (!\aluif.portOut[23]~135_combout  & (!\aluif.portOut[23]~136_combout  & ((\aluif.portOut[17]~199_combout ))))

	.dataa(\aluif.portOut[23]~135_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(\aluif.portOut[17]~197_combout ),
	.datad(\aluif.portOut[17]~199_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[17]~200_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[17]~200 .lut_mask = 16'hB9A8;
defparam \aluif.portOut[17]~200 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N16
cycloneive_lcell_comb \ShiftLeft0~98 (
// Equation(s):
// \ShiftLeft0~98_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & ((\Mux18~1_combout ))) # (!\Mux95~1_combout  & (\Mux17~1_combout ))))

	.dataa(Mux17),
	.datab(Mux18),
	.datac(Mux95),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftLeft0~98_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~98 .lut_mask = 16'hCA00;
defparam \ShiftLeft0~98 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N10
cycloneive_lcell_comb \ShiftLeft0~60 (
// Equation(s):
// \ShiftLeft0~60_combout  = (\Mux94~1_combout  & (\ShiftLeft0~49_combout )) # (!\Mux94~1_combout  & ((\ShiftLeft0~59_combout )))

	.dataa(Mux94),
	.datab(\ShiftLeft0~49_combout ),
	.datac(gnd),
	.datad(\ShiftLeft0~59_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~60_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~60 .lut_mask = 16'hDD88;
defparam \ShiftLeft0~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N30
cycloneive_lcell_comb \ShiftLeft0~106 (
// Equation(s):
// \ShiftLeft0~106_combout  = (\Mux93~2_combout  & (((\ShiftLeft0~60_combout )))) # (!\Mux93~2_combout  & ((\ShiftLeft0~99_combout ) # ((\ShiftLeft0~98_combout ))))

	.dataa(Mux931),
	.datab(\ShiftLeft0~99_combout ),
	.datac(\ShiftLeft0~98_combout ),
	.datad(\ShiftLeft0~60_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~106_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~106 .lut_mask = 16'hFE54;
defparam \ShiftLeft0~106 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N0
cycloneive_lcell_comb \ShiftLeft0~17 (
// Equation(s):
// \ShiftLeft0~17_combout  = (!\Mux92~2_combout  & (\Mux31~1_combout  & (!\Mux93~2_combout  & \ShiftLeft0~16_combout )))

	.dataa(Mux92),
	.datab(Mux31),
	.datac(Mux931),
	.datad(\ShiftLeft0~16_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~17_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~17 .lut_mask = 16'h0400;
defparam \ShiftLeft0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y25_N12
cycloneive_lcell_comb \portOut~67 (
// Equation(s):
// \portOut~67_combout  = (\Mux79~0_combout  & \Mux15~1_combout )

	.dataa(Mux79),
	.datab(gnd),
	.datac(Mux15),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~67_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~67 .lut_mask = 16'hA0A0;
defparam \portOut~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y25_N10
cycloneive_lcell_comb \aluif.portOut[16]~204 (
// Equation(s):
// \aluif.portOut[16]~204_combout  = (\aluif.portOut[15]~83_combout  & (((\portOut~67_combout ) # (!\aluif.portOut[15]~82_combout )))) # (!\aluif.portOut[15]~83_combout  & (\ShiftLeft0~17_combout  & (\aluif.portOut[15]~82_combout )))

	.dataa(\aluif.portOut[15]~83_combout ),
	.datab(\ShiftLeft0~17_combout ),
	.datac(\aluif.portOut[15]~82_combout ),
	.datad(\portOut~67_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[16]~204_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[16]~204 .lut_mask = 16'hEA4A;
defparam \aluif.portOut[16]~204 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y25_N20
cycloneive_lcell_comb \aluif.portOut[16]~205 (
// Equation(s):
// \aluif.portOut[16]~205_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[16]~204_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[16]~204_combout  & (\ShiftLeft0~43_combout )) # (!\aluif.portOut[16]~204_combout  & 
// ((\ShiftLeft0~106_combout )))))

	.dataa(\ShiftLeft0~43_combout ),
	.datab(\ShiftLeft0~106_combout ),
	.datac(\aluif.portOut[15]~81_combout ),
	.datad(\aluif.portOut[16]~204_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[16]~205_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[16]~205 .lut_mask = 16'hFA0C;
defparam \aluif.portOut[16]~205 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y25_N6
cycloneive_lcell_comb \aluif.portOut[16]~206 (
// Equation(s):
// \aluif.portOut[16]~206_combout  = (\aluif.portOut[23]~136_combout  & ((\Add0~32_combout ) # ((\aluif.portOut[23]~135_combout )))) # (!\aluif.portOut[23]~136_combout  & (((!\aluif.portOut[23]~135_combout  & \aluif.portOut[16]~205_combout ))))

	.dataa(\aluif.portOut[23]~136_combout ),
	.datab(\Add0~32_combout ),
	.datac(\aluif.portOut[23]~135_combout ),
	.datad(\aluif.portOut[16]~205_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[16]~206_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[16]~206 .lut_mask = 16'hADA8;
defparam \aluif.portOut[16]~206 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y25_N8
cycloneive_lcell_comb \portOut~68 (
// Equation(s):
// \portOut~68_combout  = \Mux79~0_combout  $ (\Mux15~1_combout )

	.dataa(Mux79),
	.datab(gnd),
	.datac(Mux15),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~68_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~68 .lut_mask = 16'h5A5A;
defparam \portOut~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N12
cycloneive_lcell_comb \portOut~66 (
// Equation(s):
// \portOut~66_combout  = (\Mux79~0_combout ) # (\Mux15~1_combout )

	.dataa(Mux79),
	.datab(gnd),
	.datac(gnd),
	.datad(Mux15),
	.cin(gnd),
	.combout(\portOut~66_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~66 .lut_mask = 16'hFFAA;
defparam \portOut~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N6
cycloneive_lcell_comb \ShiftRight0~45 (
// Equation(s):
// \ShiftRight0~45_combout  = (\ShiftRight0~41_combout ) # ((\Mux93~2_combout  & (\Mux92~2_combout  & \ShiftRight0~44_combout )))

	.dataa(\ShiftRight0~41_combout ),
	.datab(Mux931),
	.datac(Mux92),
	.datad(\ShiftRight0~44_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~45_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~45 .lut_mask = 16'hEAAA;
defparam \ShiftRight0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N26
cycloneive_lcell_comb \aluif.portOut[16]~202 (
// Equation(s):
// \aluif.portOut[16]~202_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[15]~26_combout  & \ShiftRight0~45_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~66_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(\portOut~66_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\ShiftRight0~45_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[16]~202_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[16]~202 .lut_mask = 16'hE323;
defparam \aluif.portOut[16]~202 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N4
cycloneive_lcell_comb \aluif.portOut[16]~203 (
// Equation(s):
// \aluif.portOut[16]~203_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[16]~202_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[16]~202_combout  & (!\portOut~66_combout )) # (!\aluif.portOut[16]~202_combout  & ((\Add1~32_combout )))))

	.dataa(\portOut~66_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\aluif.portOut[16]~202_combout ),
	.datad(\Add1~32_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[16]~203_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[16]~203 .lut_mask = 16'hD3D0;
defparam \aluif.portOut[16]~203 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N12
cycloneive_lcell_comb \portOut~71 (
// Equation(s):
// \portOut~71_combout  = \Mux12~1_combout  $ (\Mux76~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(Mux76),
	.cin(gnd),
	.combout(\portOut~71_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~71 .lut_mask = 16'h0FF0;
defparam \portOut~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y22_N4
cycloneive_lcell_comb \ShiftLeft0~76 (
// Equation(s):
// \ShiftLeft0~76_combout  = (!\Mux95~1_combout  & ((\Mux94~1_combout  & (\Mux14~1_combout )) # (!\Mux94~1_combout  & ((\Mux12~1_combout )))))

	.dataa(Mux95),
	.datab(Mux14),
	.datac(Mux12),
	.datad(Mux94),
	.cin(gnd),
	.combout(\ShiftLeft0~76_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~76 .lut_mask = 16'h4450;
defparam \ShiftLeft0~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N24
cycloneive_lcell_comb \ShiftLeft0~107 (
// Equation(s):
// \ShiftLeft0~107_combout  = (\Mux93~2_combout  & (\ShiftLeft0~65_combout )) # (!\Mux93~2_combout  & (((\ShiftLeft0~76_combout ) # (\ShiftLeft0~75_combout ))))

	.dataa(\ShiftLeft0~65_combout ),
	.datab(Mux931),
	.datac(\ShiftLeft0~76_combout ),
	.datad(\ShiftLeft0~75_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~107_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~107 .lut_mask = 16'hBBB8;
defparam \ShiftLeft0~107 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y22_N26
cycloneive_lcell_comb \ShiftLeft0~19 (
// Equation(s):
// \ShiftLeft0~19_combout  = (\ShiftRight0~61_combout  & ((\Mux94~1_combout  & ((\ShiftLeft0~4_combout ))) # (!\Mux94~1_combout  & (\ShiftLeft0~18_combout ))))

	.dataa(Mux94),
	.datab(\ShiftLeft0~18_combout ),
	.datac(\ShiftRight0~61_combout ),
	.datad(\ShiftLeft0~4_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~19_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~19 .lut_mask = 16'hE040;
defparam \ShiftLeft0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y22_N14
cycloneive_lcell_comb \portOut~70 (
// Equation(s):
// \portOut~70_combout  = (\Mux12~1_combout  & \Mux76~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(Mux76),
	.cin(gnd),
	.combout(\portOut~70_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~70 .lut_mask = 16'hF000;
defparam \portOut~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N8
cycloneive_lcell_comb \aluif.portOut[19]~210 (
// Equation(s):
// \aluif.portOut[19]~210_combout  = (\aluif.portOut[15]~83_combout  & (((\portOut~70_combout ) # (!\aluif.portOut[15]~82_combout )))) # (!\aluif.portOut[15]~83_combout  & (\ShiftLeft0~19_combout  & (\aluif.portOut[15]~82_combout )))

	.dataa(\aluif.portOut[15]~83_combout ),
	.datab(\ShiftLeft0~19_combout ),
	.datac(\aluif.portOut[15]~82_combout ),
	.datad(\portOut~70_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[19]~210_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[19]~210 .lut_mask = 16'hEA4A;
defparam \aluif.portOut[19]~210 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y22_N10
cycloneive_lcell_comb \aluif.portOut[19]~211 (
// Equation(s):
// \aluif.portOut[19]~211_combout  = (\aluif.portOut[15]~81_combout  & (((\aluif.portOut[19]~210_combout )))) # (!\aluif.portOut[15]~81_combout  & ((\aluif.portOut[19]~210_combout  & ((\ShiftLeft0~47_combout ))) # (!\aluif.portOut[19]~210_combout  & 
// (\ShiftLeft0~107_combout ))))

	.dataa(\aluif.portOut[15]~81_combout ),
	.datab(\ShiftLeft0~107_combout ),
	.datac(\aluif.portOut[19]~210_combout ),
	.datad(\ShiftLeft0~47_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[19]~211_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[19]~211 .lut_mask = 16'hF4A4;
defparam \aluif.portOut[19]~211 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N22
cycloneive_lcell_comb \aluif.portOut[19]~212 (
// Equation(s):
// \aluif.portOut[19]~212_combout  = (\aluif.portOut[23]~136_combout  & ((\aluif.portOut[23]~135_combout ) # ((\Add0~38_combout )))) # (!\aluif.portOut[23]~136_combout  & (!\aluif.portOut[23]~135_combout  & (\aluif.portOut[19]~211_combout )))

	.dataa(\aluif.portOut[23]~136_combout ),
	.datab(\aluif.portOut[23]~135_combout ),
	.datac(\aluif.portOut[19]~211_combout ),
	.datad(\Add0~38_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[19]~212_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[19]~212 .lut_mask = 16'hBA98;
defparam \aluif.portOut[19]~212 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N20
cycloneive_lcell_comb \portOut~69 (
// Equation(s):
// \portOut~69_combout  = (\Mux12~1_combout ) # (\Mux76~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux12),
	.datad(Mux76),
	.cin(gnd),
	.combout(\portOut~69_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~69 .lut_mask = 16'hFFF0;
defparam \portOut~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N14
cycloneive_lcell_comb \aluif.portOut[19]~208 (
// Equation(s):
// \aluif.portOut[19]~208_combout  = (\prif.ALUOP_ex [2] & (\ShiftRight0~71_combout  & ((\aluif.portOut[15]~26_combout )))) # (!\prif.ALUOP_ex [2] & (((\portOut~69_combout ) # (!\aluif.portOut[15]~26_combout ))))

	.dataa(\ShiftRight0~71_combout ),
	.datab(\portOut~69_combout ),
	.datac(prifALUOP_ex_2),
	.datad(\aluif.portOut[15]~26_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[19]~208_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[19]~208 .lut_mask = 16'hAC0F;
defparam \aluif.portOut[19]~208 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y24_N24
cycloneive_lcell_comb \aluif.portOut[19]~209 (
// Equation(s):
// \aluif.portOut[19]~209_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[19]~208_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[19]~208_combout  & ((!\portOut~69_combout ))) # (!\aluif.portOut[19]~208_combout  & (\Add1~38_combout ))))

	.dataa(prifALUOP_ex_1),
	.datab(\Add1~38_combout ),
	.datac(\aluif.portOut[19]~208_combout ),
	.datad(\portOut~69_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[19]~209_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[19]~209 .lut_mask = 16'hA4F4;
defparam \aluif.portOut[19]~209 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N26
cycloneive_lcell_comb \portOut~74 (
// Equation(s):
// \portOut~74_combout  = \Mux13~1_combout  $ (\Mux77~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux13),
	.datad(Mux77),
	.cin(gnd),
	.combout(\portOut~74_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~74 .lut_mask = 16'h0FF0;
defparam \portOut~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N10
cycloneive_lcell_comb \portOut~73 (
// Equation(s):
// \portOut~73_combout  = (\Mux13~1_combout  & \Mux77~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux13),
	.datad(Mux77),
	.cin(gnd),
	.combout(\portOut~73_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~73 .lut_mask = 16'hF000;
defparam \portOut~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N8
cycloneive_lcell_comb \aluif.portOut[18]~218 (
// Equation(s):
// \aluif.portOut[18]~218_combout  = (\aluif.portOut[15]~82_combout  & ((\aluif.portOut[15]~83_combout  & ((\portOut~73_combout ))) # (!\aluif.portOut[15]~83_combout  & (\ShiftLeft0~109_combout )))) # (!\aluif.portOut[15]~82_combout  & 
// (((\aluif.portOut[15]~83_combout ))))

	.dataa(\ShiftLeft0~109_combout ),
	.datab(\aluif.portOut[15]~82_combout ),
	.datac(\aluif.portOut[15]~83_combout ),
	.datad(\portOut~73_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[18]~218_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[18]~218 .lut_mask = 16'hF838;
defparam \aluif.portOut[18]~218 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y22_N18
cycloneive_lcell_comb \ShiftLeft0~51 (
// Equation(s):
// \ShiftLeft0~51_combout  = (\Mux93~2_combout  & ((\ShiftLeft0~35_combout ))) # (!\Mux93~2_combout  & (\ShiftLeft0~50_combout ))

	.dataa(gnd),
	.datab(\ShiftLeft0~50_combout ),
	.datac(Mux931),
	.datad(\ShiftLeft0~35_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~51_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~51 .lut_mask = 16'hFC0C;
defparam \ShiftLeft0~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N14
cycloneive_lcell_comb \aluif.portOut[18]~219 (
// Equation(s):
// \aluif.portOut[18]~219_combout  = (\aluif.portOut[18]~217_combout  & ((\aluif.portOut[15]~81_combout  & (\aluif.portOut[18]~218_combout )) # (!\aluif.portOut[15]~81_combout  & ((\ShiftLeft0~51_combout ) # (!\aluif.portOut[18]~218_combout )))))

	.dataa(\aluif.portOut[18]~217_combout ),
	.datab(\aluif.portOut[15]~81_combout ),
	.datac(\aluif.portOut[18]~218_combout ),
	.datad(\ShiftLeft0~51_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[18]~219_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[18]~219 .lut_mask = 16'hA282;
defparam \aluif.portOut[18]~219 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N28
cycloneive_lcell_comb \portOut~72 (
// Equation(s):
// \portOut~72_combout  = (\Mux13~1_combout ) # (\Mux77~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux13),
	.datad(Mux77),
	.cin(gnd),
	.combout(\portOut~72_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~72 .lut_mask = 16'hFFF0;
defparam \portOut~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N20
cycloneive_lcell_comb \aluif.portOut[18]~214 (
// Equation(s):
// \aluif.portOut[18]~214_combout  = (\prif.ALUOP_ex [2] & (\ShiftRight0~86_combout  & (\aluif.portOut[15]~26_combout ))) # (!\prif.ALUOP_ex [2] & (((\portOut~72_combout ) # (!\aluif.portOut[15]~26_combout ))))

	.dataa(\ShiftRight0~86_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\portOut~72_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[18]~214_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[18]~214 .lut_mask = 16'hB383;
defparam \aluif.portOut[18]~214 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y21_N14
cycloneive_lcell_comb \aluif.portOut[18]~215 (
// Equation(s):
// \aluif.portOut[18]~215_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[18]~214_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[18]~214_combout  & (!\portOut~72_combout )) # (!\aluif.portOut[18]~214_combout  & ((\Add1~36_combout )))))

	.dataa(prifALUOP_ex_1),
	.datab(\portOut~72_combout ),
	.datac(\Add1~36_combout ),
	.datad(\aluif.portOut[18]~214_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[18]~215_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[18]~215 .lut_mask = 16'hBB50;
defparam \aluif.portOut[18]~215 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y21_N24
cycloneive_lcell_comb \aluif.portOut[18]~220 (
// Equation(s):
// \aluif.portOut[18]~220_combout  = (\aluif.portOut[23]~135_combout  & ((\aluif.portOut[23]~136_combout ) # ((\aluif.portOut[18]~215_combout )))) # (!\aluif.portOut[23]~135_combout  & (!\aluif.portOut[23]~136_combout  & (\aluif.portOut[18]~219_combout )))

	.dataa(\aluif.portOut[23]~135_combout ),
	.datab(\aluif.portOut[23]~136_combout ),
	.datac(\aluif.portOut[18]~219_combout ),
	.datad(\aluif.portOut[18]~215_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[18]~220_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[18]~220 .lut_mask = 16'hBA98;
defparam \aluif.portOut[18]~220 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N20
cycloneive_lcell_comb \aluif.portOut[25]~226 (
// Equation(s):
// \aluif.portOut[25]~226_combout  = (\prif.ALUOP_ex [3] & ((\Mux70~0_combout  & (\prif.ALUOP_ex [0] & !\Mux6~1_combout )) # (!\Mux70~0_combout  & ((\prif.ALUOP_ex [0]) # (!\Mux6~1_combout )))))

	.dataa(Mux70),
	.datab(prifALUOP_ex_0),
	.datac(prifALUOP_ex_3),
	.datad(Mux6),
	.cin(gnd),
	.combout(\aluif.portOut[25]~226_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~226 .lut_mask = 16'h40D0;
defparam \aluif.portOut[25]~226 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N20
cycloneive_lcell_comb \ShiftLeft0~89 (
// Equation(s):
// \ShiftLeft0~89_combout  = (\Mux95~1_combout  & (\Mux94~1_combout )) # (!\Mux95~1_combout  & ((\Mux94~1_combout  & ((\Mux8~1_combout ))) # (!\Mux94~1_combout  & (\Mux6~1_combout ))))

	.dataa(Mux95),
	.datab(Mux94),
	.datac(Mux6),
	.datad(Mux8),
	.cin(gnd),
	.combout(\ShiftLeft0~89_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~89 .lut_mask = 16'hDC98;
defparam \ShiftLeft0~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N2
cycloneive_lcell_comb \ShiftLeft0~90 (
// Equation(s):
// \ShiftLeft0~90_combout  = (\ShiftLeft0~89_combout  & (((\Mux9~1_combout ) # (!\Mux95~1_combout )))) # (!\ShiftLeft0~89_combout  & (\Mux7~1_combout  & ((\Mux95~1_combout ))))

	.dataa(Mux7),
	.datab(\ShiftLeft0~89_combout ),
	.datac(Mux9),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftLeft0~90_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~90 .lut_mask = 16'hE2CC;
defparam \ShiftLeft0~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N28
cycloneive_lcell_comb \aluif.portOut[25]~222 (
// Equation(s):
// \aluif.portOut[25]~222_combout  = (\aluif.portOut[5]~52_combout  & ((\aluif.portOut[5]~51_combout ) # ((\ShiftLeft0~86_combout )))) # (!\aluif.portOut[5]~52_combout  & (!\aluif.portOut[5]~51_combout  & (\ShiftLeft0~90_combout )))

	.dataa(\aluif.portOut[5]~52_combout ),
	.datab(\aluif.portOut[5]~51_combout ),
	.datac(\ShiftLeft0~90_combout ),
	.datad(\ShiftLeft0~86_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[25]~222_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~222 .lut_mask = 16'hBA98;
defparam \aluif.portOut[25]~222 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N26
cycloneive_lcell_comb \aluif.portOut[25]~223 (
// Equation(s):
// \aluif.portOut[25]~223_combout  = (\aluif.portOut[5]~51_combout  & ((\aluif.portOut[25]~222_combout  & ((\ShiftLeft0~40_combout ))) # (!\aluif.portOut[25]~222_combout  & (\ShiftLeft0~105_combout )))) # (!\aluif.portOut[5]~51_combout  & 
// (((\aluif.portOut[25]~222_combout ))))

	.dataa(\ShiftLeft0~105_combout ),
	.datab(\aluif.portOut[5]~51_combout ),
	.datac(\ShiftLeft0~40_combout ),
	.datad(\aluif.portOut[25]~222_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[25]~223_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~223 .lut_mask = 16'hF388;
defparam \aluif.portOut[25]~223 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y23_N30
cycloneive_lcell_comb \ShiftRight0~105 (
// Equation(s):
// \ShiftRight0~105_combout  = (!\Mux92~2_combout  & ((\Mux93~2_combout  & ((\ShiftRight0~112_combout ))) # (!\Mux93~2_combout  & (\ShiftRight0~93_combout ))))

	.dataa(Mux92),
	.datab(\ShiftRight0~93_combout ),
	.datac(Mux931),
	.datad(\ShiftRight0~112_combout ),
	.cin(gnd),
	.combout(\ShiftRight0~105_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftRight0~105 .lut_mask = 16'h5404;
defparam \ShiftRight0~105 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N30
cycloneive_lcell_comb \aluif.portOut[25]~227 (
// Equation(s):
// \aluif.portOut[25]~227_combout  = (\prif.ALUOP_ex [0] & (\aluif.portOut[25]~223_combout )) # (!\prif.ALUOP_ex [0] & ((\ShiftRight0~105_combout )))

	.dataa(gnd),
	.datab(prifALUOP_ex_0),
	.datac(\aluif.portOut[25]~223_combout ),
	.datad(\ShiftRight0~105_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[25]~227_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~227 .lut_mask = 16'hF3C0;
defparam \aluif.portOut[25]~227 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y26_N22
cycloneive_lcell_comb \aluif.portOut[25]~228 (
// Equation(s):
// \aluif.portOut[25]~228_combout  = (\prif.ALUOP_ex [0] & ((\aluif.portOut[5]~55_combout ))) # (!\prif.ALUOP_ex [0] & (\aluif.portOut[15]~26_combout ))

	.dataa(gnd),
	.datab(\aluif.portOut[15]~26_combout ),
	.datac(prifALUOP_ex_0),
	.datad(\aluif.portOut[5]~55_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[25]~228_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~228 .lut_mask = 16'hFC0C;
defparam \aluif.portOut[25]~228 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N4
cycloneive_lcell_comb \aluif.portOut[25]~229 (
// Equation(s):
// \aluif.portOut[25]~229_combout  = (\prif.ALUOP_ex [2] & (((!\aluif.portOut[25]~228_combout ) # (!\aluif.portOut[25]~227_combout )))) # (!\prif.ALUOP_ex [2] & (\aluif.portOut[25]~226_combout  & ((\aluif.portOut[25]~228_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\aluif.portOut[25]~226_combout ),
	.datac(\aluif.portOut[25]~227_combout ),
	.datad(\aluif.portOut[25]~228_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[25]~229_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~229 .lut_mask = 16'h4EAA;
defparam \aluif.portOut[25]~229 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N2
cycloneive_lcell_comb \aluif.portOut[25]~225 (
// Equation(s):
// \aluif.portOut[25]~225_combout  = (\prif.ALUOP_ex [3] & ((\Mux70~0_combout  & ((\Mux6~1_combout ) # (!\prif.ALUOP_ex [0]))) # (!\Mux70~0_combout  & (\prif.ALUOP_ex [0] $ (\Mux6~1_combout )))))

	.dataa(Mux70),
	.datab(prifALUOP_ex_0),
	.datac(prifALUOP_ex_3),
	.datad(Mux6),
	.cin(gnd),
	.combout(\aluif.portOut[25]~225_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~225 .lut_mask = 16'hB060;
defparam \aluif.portOut[25]~225 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N22
cycloneive_lcell_comb \aluif.portOut[25]~230 (
// Equation(s):
// \aluif.portOut[25]~230_combout  = (\aluif.portOut[25]~225_combout  & (\prif.ALUOP_ex [1] $ (((\aluif.portOut[25]~229_combout ))))) # (!\aluif.portOut[25]~225_combout  & (\aluif.portOut[25]~226_combout  & ((!\aluif.portOut[25]~229_combout ) # 
// (!\prif.ALUOP_ex [1]))))

	.dataa(prifALUOP_ex_1),
	.datab(\aluif.portOut[25]~226_combout ),
	.datac(\aluif.portOut[25]~229_combout ),
	.datad(\aluif.portOut[25]~225_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[25]~230_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~230 .lut_mask = 16'h5A4C;
defparam \aluif.portOut[25]~230 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N22
cycloneive_lcell_comb \aluif.portOut[25]~231 (
// Equation(s):
// \aluif.portOut[25]~231_combout  = (\Mux70~0_combout ) # (\Mux6~1_combout )

	.dataa(Mux70),
	.datab(gnd),
	.datac(Mux6),
	.datad(gnd),
	.cin(gnd),
	.combout(\aluif.portOut[25]~231_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~231 .lut_mask = 16'hFAFA;
defparam \aluif.portOut[25]~231 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N8
cycloneive_lcell_comb \aluif.portOut[25]~232 (
// Equation(s):
// \aluif.portOut[25]~232_combout  = (\prif.ALUOP_ex [2] & (\ShiftRight0~105_combout  & (\aluif.portOut[15]~26_combout ))) # (!\prif.ALUOP_ex [2] & (((\aluif.portOut[25]~231_combout ) # (!\aluif.portOut[15]~26_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\ShiftRight0~105_combout ),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\aluif.portOut[25]~231_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[25]~232_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~232 .lut_mask = 16'hD585;
defparam \aluif.portOut[25]~232 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N10
cycloneive_lcell_comb \aluif.portOut[25]~233 (
// Equation(s):
// \aluif.portOut[25]~233_combout  = (\aluif.portOut[25]~230_combout  & ((\prif.ALUOP_ex [0]) # ((\aluif.portOut[25]~232_combout ) # (\Add1~50_combout ))))

	.dataa(\aluif.portOut[25]~230_combout ),
	.datab(prifALUOP_ex_0),
	.datac(\aluif.portOut[25]~232_combout ),
	.datad(\Add1~50_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[25]~233_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~233 .lut_mask = 16'hAAA8;
defparam \aluif.portOut[25]~233 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N28
cycloneive_lcell_comb \portOut~75 (
// Equation(s):
// \portOut~75_combout  = (\Mux70~0_combout  & \Mux6~1_combout )

	.dataa(Mux70),
	.datab(gnd),
	.datac(Mux6),
	.datad(gnd),
	.cin(gnd),
	.combout(\portOut~75_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~75 .lut_mask = 16'hA0A0;
defparam \portOut~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N0
cycloneive_lcell_comb \aluif.portOut[25]~224 (
// Equation(s):
// \aluif.portOut[25]~224_combout  = (\aluif.portOut[5]~55_combout  & ((\prif.ALUOP_ex [2] & (\aluif.portOut[25]~223_combout )) # (!\prif.ALUOP_ex [2] & ((\portOut~75_combout ))))) # (!\aluif.portOut[5]~55_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\aluif.portOut[25]~223_combout ),
	.datab(\portOut~75_combout ),
	.datac(\aluif.portOut[5]~55_combout ),
	.datad(prifALUOP_ex_2),
	.cin(gnd),
	.combout(\aluif.portOut[25]~224_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[25]~224 .lut_mask = 16'hA0CF;
defparam \aluif.portOut[25]~224 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N2
cycloneive_lcell_comb \portOut~77 (
// Equation(s):
// \portOut~77_combout  = (\Mux71~0_combout  & \Mux7~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux71),
	.datad(Mux7),
	.cin(gnd),
	.combout(\portOut~77_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~77 .lut_mask = 16'hF000;
defparam \portOut~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N18
cycloneive_lcell_comb \ShiftLeft0~93 (
// Equation(s):
// \ShiftLeft0~93_combout  = (\Mux94~1_combout  & ((\Mux9~1_combout ) # ((\Mux95~1_combout )))) # (!\Mux94~1_combout  & (((\Mux7~1_combout  & !\Mux95~1_combout ))))

	.dataa(Mux94),
	.datab(Mux9),
	.datac(Mux7),
	.datad(Mux95),
	.cin(gnd),
	.combout(\ShiftLeft0~93_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~93 .lut_mask = 16'hAAD8;
defparam \ShiftLeft0~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N16
cycloneive_lcell_comb \ShiftLeft0~94 (
// Equation(s):
// \ShiftLeft0~94_combout  = (\Mux95~1_combout  & ((\ShiftLeft0~93_combout  & (\Mux10~1_combout )) # (!\ShiftLeft0~93_combout  & ((\Mux8~1_combout ))))) # (!\Mux95~1_combout  & (((\ShiftLeft0~93_combout ))))

	.dataa(Mux95),
	.datab(Mux10),
	.datac(Mux8),
	.datad(\ShiftLeft0~93_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~94_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~94 .lut_mask = 16'hDDA0;
defparam \ShiftLeft0~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N18
cycloneive_lcell_comb \aluif.portOut[24]~235 (
// Equation(s):
// \aluif.portOut[24]~235_combout  = (\aluif.portOut[5]~51_combout  & ((\aluif.portOut[5]~52_combout ) # ((\ShiftLeft0~106_combout )))) # (!\aluif.portOut[5]~51_combout  & (!\aluif.portOut[5]~52_combout  & ((\ShiftLeft0~94_combout ))))

	.dataa(\aluif.portOut[5]~51_combout ),
	.datab(\aluif.portOut[5]~52_combout ),
	.datac(\ShiftLeft0~106_combout ),
	.datad(\ShiftLeft0~94_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[24]~235_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[24]~235 .lut_mask = 16'hB9A8;
defparam \aluif.portOut[24]~235 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N20
cycloneive_lcell_comb \aluif.portOut[24]~236 (
// Equation(s):
// \aluif.portOut[24]~236_combout  = (\aluif.portOut[5]~52_combout  & ((\aluif.portOut[24]~235_combout  & (\ShiftLeft0~44_combout )) # (!\aluif.portOut[24]~235_combout  & ((\ShiftLeft0~97_combout ))))) # (!\aluif.portOut[5]~52_combout  & 
// (((\aluif.portOut[24]~235_combout ))))

	.dataa(\ShiftLeft0~44_combout ),
	.datab(\aluif.portOut[5]~52_combout ),
	.datac(\ShiftLeft0~97_combout ),
	.datad(\aluif.portOut[24]~235_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[24]~236_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[24]~236 .lut_mask = 16'hBBC0;
defparam \aluif.portOut[24]~236 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N12
cycloneive_lcell_comb \aluif.portOut[24]~237 (
// Equation(s):
// \aluif.portOut[24]~237_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[5]~55_combout  & \aluif.portOut[24]~236_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~77_combout ) # ((!\aluif.portOut[5]~55_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\portOut~77_combout ),
	.datac(\aluif.portOut[5]~55_combout ),
	.datad(\aluif.portOut[24]~236_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[24]~237_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[24]~237 .lut_mask = 16'hE545;
defparam \aluif.portOut[24]~237 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N24
cycloneive_lcell_comb \portOut~76 (
// Equation(s):
// \portOut~76_combout  = \Mux71~0_combout  $ (\Mux7~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux71),
	.datad(Mux7),
	.cin(gnd),
	.combout(\portOut~76_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~76 .lut_mask = 16'h0FF0;
defparam \portOut~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y21_N30
cycloneive_lcell_comb \aluif.portOut[24]~238 (
// Equation(s):
// \aluif.portOut[24]~238_combout  = (\aluif.portOut[24]~237_combout  & ((\prif.ALUOP_ex [1]) # ((\portOut~76_combout )))) # (!\aluif.portOut[24]~237_combout  & (!\prif.ALUOP_ex [1] & (\Add0~48_combout )))

	.dataa(\aluif.portOut[24]~237_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\Add0~48_combout ),
	.datad(\portOut~76_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[24]~238_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[24]~238 .lut_mask = 16'hBA98;
defparam \aluif.portOut[24]~238 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N10
cycloneive_lcell_comb \portOut~78 (
// Equation(s):
// \portOut~78_combout  = (\Mux7~1_combout ) # (\Mux71~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux7),
	.datad(Mux71),
	.cin(gnd),
	.combout(\portOut~78_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~78 .lut_mask = 16'hFFF0;
defparam \portOut~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N28
cycloneive_lcell_comb \aluif.portOut[24]~239 (
// Equation(s):
// \aluif.portOut[24]~239_combout  = (\prif.ALUOP_ex [2] & (((\aluif.portOut[15]~26_combout  & \ShiftRight0~106_combout )))) # (!\prif.ALUOP_ex [2] & ((\portOut~78_combout ) # ((!\aluif.portOut[15]~26_combout ))))

	.dataa(\portOut~78_combout ),
	.datab(prifALUOP_ex_2),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\ShiftRight0~106_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[24]~239_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[24]~239 .lut_mask = 16'hE323;
defparam \aluif.portOut[24]~239 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y23_N14
cycloneive_lcell_comb \aluif.portOut[24]~240 (
// Equation(s):
// \aluif.portOut[24]~240_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[24]~239_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[24]~239_combout  & (!\portOut~78_combout )) # (!\aluif.portOut[24]~239_combout  & ((\Add1~48_combout )))))

	.dataa(\portOut~78_combout ),
	.datab(prifALUOP_ex_1),
	.datac(\Add1~48_combout ),
	.datad(\aluif.portOut[24]~239_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[24]~240_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[24]~240 .lut_mask = 16'hDD30;
defparam \aluif.portOut[24]~240 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N16
cycloneive_lcell_comb \portOut~80 (
// Equation(s):
// \portOut~80_combout  = (\Mux4~1_combout ) # (\Mux68~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux4),
	.datad(Mux68),
	.cin(gnd),
	.combout(\portOut~80_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~80 .lut_mask = 16'hFFF0;
defparam \portOut~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N6
cycloneive_lcell_comb \aluif.portOut[27]~247 (
// Equation(s):
// \aluif.portOut[27]~247_combout  = (\aluif.portOut[15]~26_combout  & ((\prif.ALUOP_ex [2] & ((\ShiftRight0~107_combout ))) # (!\prif.ALUOP_ex [2] & (\portOut~80_combout )))) # (!\aluif.portOut[15]~26_combout  & (((!\prif.ALUOP_ex [2]))))

	.dataa(\aluif.portOut[15]~26_combout ),
	.datab(\portOut~80_combout ),
	.datac(prifALUOP_ex_2),
	.datad(\ShiftRight0~107_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[27]~247_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[27]~247 .lut_mask = 16'hAD0D;
defparam \aluif.portOut[27]~247 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N20
cycloneive_lcell_comb \aluif.portOut[27]~248 (
// Equation(s):
// \aluif.portOut[27]~248_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[27]~247_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[27]~247_combout  & (!\portOut~80_combout )) # (!\aluif.portOut[27]~247_combout  & ((\Add1~54_combout )))))

	.dataa(prifALUOP_ex_1),
	.datab(\portOut~80_combout ),
	.datac(\Add1~54_combout ),
	.datad(\aluif.portOut[27]~247_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[27]~248_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[27]~248 .lut_mask = 16'hBB50;
defparam \aluif.portOut[27]~248 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N4
cycloneive_lcell_comb \aluif.portOut[27]~245 (
// Equation(s):
// \aluif.portOut[27]~245_combout  = \Mux4~1_combout  $ (\Mux68~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux4),
	.datad(Mux68),
	.cin(gnd),
	.combout(\aluif.portOut[27]~245_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[27]~245 .lut_mask = 16'h0FF0;
defparam \aluif.portOut[27]~245 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N24
cycloneive_lcell_comb \portOut~79 (
// Equation(s):
// \portOut~79_combout  = (\Mux4~1_combout  & \Mux68~0_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux4),
	.datad(Mux68),
	.cin(gnd),
	.combout(\portOut~79_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~79 .lut_mask = 16'hF000;
defparam \portOut~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N10
cycloneive_lcell_comb \aluif.portOut[27]~244 (
// Equation(s):
// \aluif.portOut[27]~244_combout  = (\prif.ALUOP_ex [2] & (\aluif.portOut[27]~243_combout  & ((\aluif.portOut[5]~55_combout )))) # (!\prif.ALUOP_ex [2] & (((\portOut~79_combout ) # (!\aluif.portOut[5]~55_combout ))))

	.dataa(\aluif.portOut[27]~243_combout ),
	.datab(\portOut~79_combout ),
	.datac(prifALUOP_ex_2),
	.datad(\aluif.portOut[5]~55_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[27]~244_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[27]~244 .lut_mask = 16'hAC0F;
defparam \aluif.portOut[27]~244 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y24_N18
cycloneive_lcell_comb \aluif.portOut[27]~246 (
// Equation(s):
// \aluif.portOut[27]~246_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[27]~244_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[27]~244_combout  & ((\aluif.portOut[27]~245_combout ))) # (!\aluif.portOut[27]~244_combout  & (\Add0~54_combout ))))

	.dataa(prifALUOP_ex_1),
	.datab(\Add0~54_combout ),
	.datac(\aluif.portOut[27]~245_combout ),
	.datad(\aluif.portOut[27]~244_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[27]~246_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[27]~246 .lut_mask = 16'hFA44;
defparam \aluif.portOut[27]~246 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y23_N30
cycloneive_lcell_comb \portOut~82 (
// Equation(s):
// \portOut~82_combout  = (\Mux69~0_combout ) # (\Mux5~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux69),
	.datad(Mux5),
	.cin(gnd),
	.combout(\portOut~82_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~82 .lut_mask = 16'hFFF0;
defparam \portOut~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N18
cycloneive_lcell_comb \aluif.portOut[26]~255 (
// Equation(s):
// \aluif.portOut[26]~255_combout  = (\prif.ALUOP_ex [2] & (\ShiftRight0~108_combout  & (\aluif.portOut[15]~26_combout ))) # (!\prif.ALUOP_ex [2] & (((\portOut~82_combout ) # (!\aluif.portOut[15]~26_combout ))))

	.dataa(prifALUOP_ex_2),
	.datab(\ShiftRight0~108_combout ),
	.datac(\aluif.portOut[15]~26_combout ),
	.datad(\portOut~82_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[26]~255_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[26]~255 .lut_mask = 16'hD585;
defparam \aluif.portOut[26]~255 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N12
cycloneive_lcell_comb \aluif.portOut[26]~256 (
// Equation(s):
// \aluif.portOut[26]~256_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[26]~255_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[26]~255_combout  & (!\portOut~82_combout )) # (!\aluif.portOut[26]~255_combout  & ((\Add1~52_combout )))))

	.dataa(\portOut~82_combout ),
	.datab(\Add1~52_combout ),
	.datac(prifALUOP_ex_1),
	.datad(\aluif.portOut[26]~255_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[26]~256_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[26]~256 .lut_mask = 16'hF50C;
defparam \aluif.portOut[26]~256 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y23_N12
cycloneive_lcell_comb \aluif.portOut[26]~253 (
// Equation(s):
// \aluif.portOut[26]~253_combout  = \Mux69~0_combout  $ (\Mux5~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux69),
	.datad(Mux5),
	.cin(gnd),
	.combout(\aluif.portOut[26]~253_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[26]~253 .lut_mask = 16'h0FF0;
defparam \aluif.portOut[26]~253 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y23_N30
cycloneive_lcell_comb \portOut~81 (
// Equation(s):
// \portOut~81_combout  = (\Mux69~0_combout  & \Mux5~1_combout )

	.dataa(gnd),
	.datab(gnd),
	.datac(Mux69),
	.datad(Mux5),
	.cin(gnd),
	.combout(\portOut~81_combout ),
	.cout());
// synopsys translate_off
defparam \portOut~81 .lut_mask = 16'hF000;
defparam \portOut~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N4
cycloneive_lcell_comb \ShiftLeft0~103 (
// Equation(s):
// \ShiftLeft0~103_combout  = (\Mux94~1_combout  & ((\Mux95~1_combout  & (\Mux8~1_combout )) # (!\Mux95~1_combout  & ((\Mux7~1_combout )))))

	.dataa(Mux94),
	.datab(Mux95),
	.datac(Mux8),
	.datad(Mux7),
	.cin(gnd),
	.combout(\ShiftLeft0~103_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~103 .lut_mask = 16'hA280;
defparam \ShiftLeft0~103 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y23_N30
cycloneive_lcell_comb \ShiftLeft0~104 (
// Equation(s):
// \ShiftLeft0~104_combout  = (\ShiftLeft0~103_combout ) # ((!\Mux94~1_combout  & \ShiftLeft0~92_combout ))

	.dataa(gnd),
	.datab(Mux94),
	.datac(\ShiftLeft0~103_combout ),
	.datad(\ShiftLeft0~92_combout ),
	.cin(gnd),
	.combout(\ShiftLeft0~104_combout ),
	.cout());
// synopsys translate_off
defparam \ShiftLeft0~104 .lut_mask = 16'hF3F0;
defparam \ShiftLeft0~104 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N12
cycloneive_lcell_comb \aluif.portOut[26]~250 (
// Equation(s):
// \aluif.portOut[26]~250_combout  = (\aluif.portOut[5]~52_combout  & (((\aluif.portOut[5]~51_combout )))) # (!\aluif.portOut[5]~52_combout  & ((\aluif.portOut[5]~51_combout  & (\ShiftLeft0~108_combout )) # (!\aluif.portOut[5]~51_combout  & 
// ((\ShiftLeft0~104_combout )))))

	.dataa(\ShiftLeft0~108_combout ),
	.datab(\aluif.portOut[5]~52_combout ),
	.datac(\aluif.portOut[5]~51_combout ),
	.datad(\ShiftLeft0~104_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[26]~250_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[26]~250 .lut_mask = 16'hE3E0;
defparam \aluif.portOut[26]~250 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y22_N10
cycloneive_lcell_comb \aluif.portOut[26]~251 (
// Equation(s):
// \aluif.portOut[26]~251_combout  = (\aluif.portOut[5]~52_combout  & ((\aluif.portOut[26]~250_combout  & (\ShiftLeft0~52_combout )) # (!\aluif.portOut[26]~250_combout  & ((\ShiftLeft0~79_combout ))))) # (!\aluif.portOut[5]~52_combout  & 
// (((\aluif.portOut[26]~250_combout ))))

	.dataa(\ShiftLeft0~52_combout ),
	.datab(\aluif.portOut[5]~52_combout ),
	.datac(\ShiftLeft0~79_combout ),
	.datad(\aluif.portOut[26]~250_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[26]~251_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[26]~251 .lut_mask = 16'hBBC0;
defparam \aluif.portOut[26]~251 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N6
cycloneive_lcell_comb \aluif.portOut[26]~252 (
// Equation(s):
// \aluif.portOut[26]~252_combout  = (\prif.ALUOP_ex [2] & (\aluif.portOut[5]~55_combout  & ((\aluif.portOut[26]~251_combout )))) # (!\prif.ALUOP_ex [2] & (((\portOut~81_combout )) # (!\aluif.portOut[5]~55_combout )))

	.dataa(prifALUOP_ex_2),
	.datab(\aluif.portOut[5]~55_combout ),
	.datac(\portOut~81_combout ),
	.datad(\aluif.portOut[26]~251_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[26]~252_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[26]~252 .lut_mask = 16'hD951;
defparam \aluif.portOut[26]~252 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y22_N16
cycloneive_lcell_comb \aluif.portOut[26]~254 (
// Equation(s):
// \aluif.portOut[26]~254_combout  = (\prif.ALUOP_ex [1] & (((\aluif.portOut[26]~252_combout )))) # (!\prif.ALUOP_ex [1] & ((\aluif.portOut[26]~252_combout  & ((\aluif.portOut[26]~253_combout ))) # (!\aluif.portOut[26]~252_combout  & (\Add0~52_combout ))))

	.dataa(prifALUOP_ex_1),
	.datab(\Add0~52_combout ),
	.datac(\aluif.portOut[26]~253_combout ),
	.datad(\aluif.portOut[26]~252_combout ),
	.cin(gnd),
	.combout(\aluif.portOut[26]~254_combout ),
	.cout());
// synopsys translate_off
defparam \aluif.portOut[26]~254 .lut_mask = 16'hFA44;
defparam \aluif.portOut[26]~254 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module control_unit (
	prifimemload_id_31,
	prifimemload_id_30,
	prifimemload_id_29,
	prifimemload_id_27,
	prifimemload_id_26,
	prifimemload_id_28,
	prifimemload_id_3,
	prifimemload_id_1,
	prifimemload_id_5,
	prifimemload_id_4,
	prifimemload_id_2,
	prifimemload_id_0,
	Equal15,
	Equal11,
	Equal0,
	Equal10,
	Equal12,
	Equal20,
	Equal26,
	Equal25,
	Equal13,
	dataScr_ex,
	WideNor0,
	Selector0,
	Equal4,
	Selector2,
	Selector21,
	ALUScr_ex,
	Selector3,
	Equal131,
	ALUScr_ex1,
	devpor,
	devclrn,
	devoe);
input 	prifimemload_id_31;
input 	prifimemload_id_30;
input 	prifimemload_id_29;
input 	prifimemload_id_27;
input 	prifimemload_id_26;
input 	prifimemload_id_28;
input 	prifimemload_id_3;
input 	prifimemload_id_1;
input 	prifimemload_id_5;
input 	prifimemload_id_4;
input 	prifimemload_id_2;
input 	prifimemload_id_0;
output 	Equal15;
output 	Equal11;
output 	Equal0;
output 	Equal10;
output 	Equal12;
output 	Equal20;
output 	Equal26;
output 	Equal25;
output 	Equal13;
input 	dataScr_ex;
output 	WideNor0;
output 	Selector0;
output 	Equal4;
output 	Selector2;
output 	Selector21;
input 	ALUScr_ex;
output 	Selector3;
output 	Equal131;
input 	ALUScr_ex1;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Equal25~0_combout ;
wire \Equal16~0_combout ;
wire \WideNor0~0_combout ;
wire \WideNor0~1_combout ;
wire \Selector3~0_combout ;
wire \Selector0~0_combout ;
wire \Selector0~1_combout ;
wire \Selector2~6_combout ;
wire \Selector2~7_combout ;
wire \Selector3~2_combout ;
wire \Selector3~3_combout ;
wire \Selector3~4_combout ;
wire \Selector3~1_combout ;


// Location: LCCOMB_X53_Y31_N28
cycloneive_lcell_comb \Equal15~0 (
// Equation(s):
// Equal15 = (!\prif.imemload_id [30] & (!\prif.imemload_id [29] & (!\prif.imemload_id [27] & !\prif.imemload_id [31])))

	.dataa(prifimemload_id_30),
	.datab(prifimemload_id_29),
	.datac(prifimemload_id_27),
	.datad(prifimemload_id_31),
	.cin(gnd),
	.combout(Equal15),
	.cout());
// synopsys translate_off
defparam \Equal15~0 .lut_mask = 16'h0001;
defparam \Equal15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N26
cycloneive_lcell_comb \Equal11~0 (
// Equation(s):
// Equal11 = (!\prif.imemload_id [26] & (Equal15 & !\prif.imemload_id [28]))

	.dataa(gnd),
	.datab(prifimemload_id_26),
	.datac(Equal15),
	.datad(prifimemload_id_28),
	.cin(gnd),
	.combout(Equal11),
	.cout());
// synopsys translate_off
defparam \Equal11~0 .lut_mask = 16'h0030;
defparam \Equal11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N18
cycloneive_lcell_comb \Equal0~0 (
// Equation(s):
// Equal0 = (!\prif.imemload_id [5] & (!\prif.imemload_id [4] & (!\prif.imemload_id [2] & !\prif.imemload_id [0])))

	.dataa(prifimemload_id_5),
	.datab(prifimemload_id_4),
	.datac(prifimemload_id_2),
	.datad(prifimemload_id_0),
	.cin(gnd),
	.combout(Equal0),
	.cout());
// synopsys translate_off
defparam \Equal0~0 .lut_mask = 16'h0001;
defparam \Equal0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N20
cycloneive_lcell_comb \Equal10~0 (
// Equation(s):
// Equal10 = ((\prif.imemload_id [1]) # (!Equal0)) # (!\prif.imemload_id [3])

	.dataa(gnd),
	.datab(prifimemload_id_3),
	.datac(Equal0),
	.datad(prifimemload_id_1),
	.cin(gnd),
	.combout(Equal10),
	.cout());
// synopsys translate_off
defparam \Equal10~0 .lut_mask = 16'hFF3F;
defparam \Equal10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N18
cycloneive_lcell_comb \Equal12~0 (
// Equation(s):
// Equal12 = (\prif.imemload_id [27] & (!\prif.imemload_id [30] & (!\prif.imemload_id [29] & !\prif.imemload_id [28])))

	.dataa(prifimemload_id_27),
	.datab(prifimemload_id_30),
	.datac(prifimemload_id_29),
	.datad(prifimemload_id_28),
	.cin(gnd),
	.combout(Equal12),
	.cout());
// synopsys translate_off
defparam \Equal12~0 .lut_mask = 16'h0002;
defparam \Equal12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N0
cycloneive_lcell_comb \Equal20~0 (
// Equation(s):
// Equal20 = (\prif.imemload_id [29] & (!\prif.imemload_id [30] & (!\prif.imemload_id [31] & \prif.imemload_id [28])))

	.dataa(prifimemload_id_29),
	.datab(prifimemload_id_30),
	.datac(prifimemload_id_31),
	.datad(prifimemload_id_28),
	.cin(gnd),
	.combout(Equal20),
	.cout());
// synopsys translate_off
defparam \Equal20~0 .lut_mask = 16'h0200;
defparam \Equal20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N28
cycloneive_lcell_comb \Equal26~0 (
// Equation(s):
// Equal26 = (\prif.imemload_id [28] & (\Equal25~0_combout  & \prif.imemload_id [30]))

	.dataa(prifimemload_id_28),
	.datab(gnd),
	.datac(\Equal25~0_combout ),
	.datad(prifimemload_id_30),
	.cin(gnd),
	.combout(Equal26),
	.cout());
// synopsys translate_off
defparam \Equal26~0 .lut_mask = 16'hA000;
defparam \Equal26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N28
cycloneive_lcell_comb \Equal25~1 (
// Equation(s):
// Equal25 = (\Equal25~0_combout  & (!\prif.imemload_id [30] & !\prif.imemload_id [28]))

	.dataa(\Equal25~0_combout ),
	.datab(prifimemload_id_30),
	.datac(gnd),
	.datad(prifimemload_id_28),
	.cin(gnd),
	.combout(Equal25),
	.cout());
// synopsys translate_off
defparam \Equal25~1 .lut_mask = 16'h0022;
defparam \Equal25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N10
cycloneive_lcell_comb \Equal13~0 (
// Equation(s):
// Equal13 = (\prif.imemload_id [26] & (!\prif.imemload_id [31] & Equal12))

	.dataa(prifimemload_id_26),
	.datab(gnd),
	.datac(prifimemload_id_31),
	.datad(Equal12),
	.cin(gnd),
	.combout(Equal13),
	.cout());
// synopsys translate_off
defparam \Equal13~0 .lut_mask = 16'h0A00;
defparam \Equal13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N2
cycloneive_lcell_comb \WideNor0~2 (
// Equation(s):
// WideNor0 = (\WideNor0~1_combout  & (dataScr_ex & ((\prif.imemload_id [27]) # (!Equal20))))

	.dataa(\WideNor0~1_combout ),
	.datab(prifimemload_id_27),
	.datac(Equal20),
	.datad(dataScr_ex),
	.cin(gnd),
	.combout(WideNor0),
	.cout());
// synopsys translate_off
defparam \WideNor0~2 .lut_mask = 16'h8A00;
defparam \WideNor0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N14
cycloneive_lcell_comb \Selector0~2 (
// Equation(s):
// Selector0 = (((Equal11 & \Selector0~0_combout )) # (!ALUScr_ex3)) # (!\Selector0~1_combout )

	.dataa(Equal11),
	.datab(\Selector0~0_combout ),
	.datac(\Selector0~1_combout ),
	.datad(ALUScr_ex1),
	.cin(gnd),
	.combout(Selector0),
	.cout());
// synopsys translate_off
defparam \Selector0~2 .lut_mask = 16'h8FFF;
defparam \Selector0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N30
cycloneive_lcell_comb \Equal4~0 (
// Equation(s):
// Equal4 = (\prif.imemload_id [5] & (!\prif.imemload_id [3] & (\prif.imemload_id [2] & !\prif.imemload_id [4])))

	.dataa(prifimemload_id_5),
	.datab(prifimemload_id_3),
	.datac(prifimemload_id_2),
	.datad(prifimemload_id_4),
	.cin(gnd),
	.combout(Equal4),
	.cout());
// synopsys translate_off
defparam \Equal4~0 .lut_mask = 16'h0020;
defparam \Equal4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N0
cycloneive_lcell_comb \Selector2~4 (
// Equation(s):
// Selector2 = (Equal10 & (!\prif.imemload_id [26] & (Equal15 & !\prif.imemload_id [28])))

	.dataa(Equal10),
	.datab(prifimemload_id_26),
	.datac(Equal15),
	.datad(prifimemload_id_28),
	.cin(gnd),
	.combout(Selector2),
	.cout());
// synopsys translate_off
defparam \Selector2~4 .lut_mask = 16'h0020;
defparam \Selector2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N20
cycloneive_lcell_comb \Selector2~5 (
// Equation(s):
// Selector21 = (\Selector2~6_combout ) # (((Selector2 & \Selector2~7_combout )) # (!\WideNor0~1_combout ))

	.dataa(\Selector2~6_combout ),
	.datab(Selector2),
	.datac(\Selector2~7_combout ),
	.datad(\WideNor0~1_combout ),
	.cin(gnd),
	.combout(Selector21),
	.cout());
// synopsys translate_off
defparam \Selector2~5 .lut_mask = 16'hEAFF;
defparam \Selector2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N24
cycloneive_lcell_comb \Selector3~5 (
// Equation(s):
// Selector3 = (\Selector3~1_combout ) # (((Equal11 & \Selector3~4_combout )) # (!ALUScr_ex2))

	.dataa(Equal11),
	.datab(\Selector3~4_combout ),
	.datac(\Selector3~1_combout ),
	.datad(ALUScr_ex),
	.cin(gnd),
	.combout(Selector3),
	.cout());
// synopsys translate_off
defparam \Selector3~5 .lut_mask = 16'hF8FF;
defparam \Selector3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N2
cycloneive_lcell_comb \Equal13~1 (
// Equation(s):
// Equal131 = (\prif.imemload_id [26] & Equal12)

	.dataa(gnd),
	.datab(prifimemload_id_26),
	.datac(gnd),
	.datad(Equal12),
	.cin(gnd),
	.combout(Equal131),
	.cout());
// synopsys translate_off
defparam \Equal13~1 .lut_mask = 16'hCC00;
defparam \Equal13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N6
cycloneive_lcell_comb \Equal25~0 (
// Equation(s):
// \Equal25~0_combout  = (\prif.imemload_id [27] & (\prif.imemload_id [31] & (\prif.imemload_id [29] & \prif.imemload_id [26])))

	.dataa(prifimemload_id_27),
	.datab(prifimemload_id_31),
	.datac(prifimemload_id_29),
	.datad(prifimemload_id_26),
	.cin(gnd),
	.combout(\Equal25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal25~0 .lut_mask = 16'h8000;
defparam \Equal25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N8
cycloneive_lcell_comb \Equal16~0 (
// Equation(s):
// \Equal16~0_combout  = (\prif.imemload_id [29] & (!\prif.imemload_id [30] & (!\prif.imemload_id [31] & !\prif.imemload_id [28])))

	.dataa(prifimemload_id_29),
	.datab(prifimemload_id_30),
	.datac(prifimemload_id_31),
	.datad(prifimemload_id_28),
	.cin(gnd),
	.combout(\Equal16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal16~0 .lut_mask = 16'h0002;
defparam \Equal16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N26
cycloneive_lcell_comb \WideNor0~0 (
// Equation(s):
// \WideNor0~0_combout  = (!\Equal16~0_combout  & (((\prif.imemload_id [26]) # (!Equal20)) # (!\prif.imemload_id [27])))

	.dataa(prifimemload_id_27),
	.datab(Equal20),
	.datac(\Equal16~0_combout ),
	.datad(prifimemload_id_26),
	.cin(gnd),
	.combout(\WideNor0~0_combout ),
	.cout());
// synopsys translate_off
defparam \WideNor0~0 .lut_mask = 16'h0F07;
defparam \WideNor0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N16
cycloneive_lcell_comb \WideNor0~1 (
// Equation(s):
// \WideNor0~1_combout  = (\WideNor0~0_combout  & (((!\prif.imemload_id [26]) # (!\prif.imemload_id [31])) # (!Equal12)))

	.dataa(Equal12),
	.datab(prifimemload_id_31),
	.datac(\WideNor0~0_combout ),
	.datad(prifimemload_id_26),
	.cin(gnd),
	.combout(\WideNor0~1_combout ),
	.cout());
// synopsys translate_off
defparam \WideNor0~1 .lut_mask = 16'h70F0;
defparam \WideNor0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N4
cycloneive_lcell_comb \Selector3~0 (
// Equation(s):
// \Selector3~0_combout  = (!\prif.imemload_id [4] & (\prif.imemload_id [5] & \prif.imemload_id [1]))

	.dataa(gnd),
	.datab(prifimemload_id_4),
	.datac(prifimemload_id_5),
	.datad(prifimemload_id_1),
	.cin(gnd),
	.combout(\Selector3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~0 .lut_mask = 16'h3000;
defparam \Selector3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N20
cycloneive_lcell_comb \Selector0~0 (
// Equation(s):
// \Selector0~0_combout  = ((!\prif.imemload_id [2] & (\Selector3~0_combout  & \prif.imemload_id [3]))) # (!Equal10)

	.dataa(Equal10),
	.datab(prifimemload_id_2),
	.datac(\Selector3~0_combout ),
	.datad(prifimemload_id_3),
	.cin(gnd),
	.combout(\Selector0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~0 .lut_mask = 16'h7555;
defparam \Selector0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N22
cycloneive_lcell_comb \Selector0~1 (
// Equation(s):
// \Selector0~1_combout  = (!\prif.imemload_id [27]) # (!\Equal16~0_combout )

	.dataa(gnd),
	.datab(\Equal16~0_combout ),
	.datac(gnd),
	.datad(prifimemload_id_27),
	.cin(gnd),
	.combout(\Selector0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector0~1 .lut_mask = 16'h33FF;
defparam \Selector0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N12
cycloneive_lcell_comb \Selector2~6 (
// Equation(s):
// \Selector2~6_combout  = (\prif.imemload_id [28] & (((Equal15)))) # (!\prif.imemload_id [28] & (\Equal25~0_combout  & (!\prif.imemload_id [30])))

	.dataa(\Equal25~0_combout ),
	.datab(prifimemload_id_30),
	.datac(Equal15),
	.datad(prifimemload_id_28),
	.cin(gnd),
	.combout(\Selector2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~6 .lut_mask = 16'hF022;
defparam \Selector2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N2
cycloneive_lcell_comb \Selector2~7 (
// Equation(s):
// \Selector2~7_combout  = (\prif.imemload_id [3] & (((\prif.imemload_id [1]) # (!Equal4)))) # (!\prif.imemload_id [3] & (!Equal0 & ((\prif.imemload_id [1]) # (!Equal4))))

	.dataa(prifimemload_id_3),
	.datab(Equal0),
	.datac(Equal4),
	.datad(prifimemload_id_1),
	.cin(gnd),
	.combout(\Selector2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Selector2~7 .lut_mask = 16'hBB0B;
defparam \Selector2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N8
cycloneive_lcell_comb \Selector3~2 (
// Equation(s):
// \Selector3~2_combout  = (\Selector3~0_combout  & ((\prif.imemload_id [3] & (!\prif.imemload_id [2] & \prif.imemload_id [0])) # (!\prif.imemload_id [3] & ((\prif.imemload_id [0]) # (!\prif.imemload_id [2])))))

	.dataa(\Selector3~0_combout ),
	.datab(prifimemload_id_3),
	.datac(prifimemload_id_2),
	.datad(prifimemload_id_0),
	.cin(gnd),
	.combout(\Selector3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~2 .lut_mask = 16'h2A02;
defparam \Selector3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N10
cycloneive_lcell_comb \Selector3~3 (
// Equation(s):
// \Selector3~3_combout  = (\Selector3~2_combout ) # ((!\prif.imemload_id [3] & (Equal0 & \prif.imemload_id [1])))

	.dataa(prifimemload_id_3),
	.datab(Equal0),
	.datac(\Selector3~2_combout ),
	.datad(prifimemload_id_1),
	.cin(gnd),
	.combout(\Selector3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~3 .lut_mask = 16'hF4F0;
defparam \Selector3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N12
cycloneive_lcell_comb \Selector3~4 (
// Equation(s):
// \Selector3~4_combout  = (\Selector3~3_combout ) # ((\prif.imemload_id [0] & (Equal4 & !\prif.imemload_id [1])))

	.dataa(\Selector3~3_combout ),
	.datab(prifimemload_id_0),
	.datac(Equal4),
	.datad(prifimemload_id_1),
	.cin(gnd),
	.combout(\Selector3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~4 .lut_mask = 16'hAAEA;
defparam \Selector3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N10
cycloneive_lcell_comb \Selector3~1 (
// Equation(s):
// \Selector3~1_combout  = (\prif.imemload_id [26] & ((\prif.imemload_id [27] & ((\Equal16~0_combout ))) # (!\prif.imemload_id [27] & (Equal20))))

	.dataa(prifimemload_id_27),
	.datab(Equal20),
	.datac(\Equal16~0_combout ),
	.datad(prifimemload_id_26),
	.cin(gnd),
	.combout(\Selector3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Selector3~1 .lut_mask = 16'hE400;
defparam \Selector3~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module hazard_unit (
	prifRegwen_mem,
	prifregwrite_mem_4,
	prifregwrite_mem_0,
	prifregwrite_mem_1,
	prifregwrite_mem_2,
	prifregwrite_mem_3,
	prifrt_ex_1,
	prifrt_ex_0,
	prifrt_ex_3,
	prifrt_ex_2,
	prifrt_ex_4,
	prifopcode_mem_1,
	prifopcode_mem_0,
	prifopcode_mem_2,
	prifopcode_mem_3,
	prifopcode_mem_5,
	prifopcode_mem_4,
	prifzero_flag_mem,
	prifinstr_mem_3,
	prifinstr_mem_5,
	prifinstr_mem_4,
	prifinstr_mem_2,
	prifinstr_mem_1,
	prifinstr_mem_0,
	prifopcode_ex_5,
	prifopcode_ex_0,
	prifopcode_ex_1,
	prifopcode_ex_2,
	prifopcode_ex_4,
	LessThan1,
	always0,
	ptBScr,
	prifRegwen_wb,
	prifregwrite_wb_2,
	prifregwrite_wb_0,
	prifregwrite_wb_1,
	prifregwrite_wb_4,
	prifregwrite_wb_3,
	Equal8,
	always01,
	prifrs_ex_1,
	prifrs_ex_0,
	prifrs_ex_3,
	prifrs_ex_2,
	prifrs_ex_4,
	always02,
	ptAScr,
	always03,
	exmem_en,
	Equal1,
	ccifiwait_0,
	always1,
	ifid_en,
	pc_en,
	flush_idex,
	prifhalt_wb,
	ifid_en1,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	prifRegwen_mem;
input 	prifregwrite_mem_4;
input 	prifregwrite_mem_0;
input 	prifregwrite_mem_1;
input 	prifregwrite_mem_2;
input 	prifregwrite_mem_3;
input 	prifrt_ex_1;
input 	prifrt_ex_0;
input 	prifrt_ex_3;
input 	prifrt_ex_2;
input 	prifrt_ex_4;
input 	prifopcode_mem_1;
input 	prifopcode_mem_0;
input 	prifopcode_mem_2;
input 	prifopcode_mem_3;
input 	prifopcode_mem_5;
input 	prifopcode_mem_4;
input 	prifzero_flag_mem;
input 	prifinstr_mem_3;
input 	prifinstr_mem_5;
input 	prifinstr_mem_4;
input 	prifinstr_mem_2;
input 	prifinstr_mem_1;
input 	prifinstr_mem_0;
input 	prifopcode_ex_5;
input 	prifopcode_ex_0;
input 	prifopcode_ex_1;
input 	prifopcode_ex_2;
input 	prifopcode_ex_4;
input 	LessThan1;
input 	always0;
output 	ptBScr;
input 	prifRegwen_wb;
input 	prifregwrite_wb_2;
input 	prifregwrite_wb_0;
input 	prifregwrite_wb_1;
input 	prifregwrite_wb_4;
input 	prifregwrite_wb_3;
output 	Equal8;
output 	always01;
input 	prifrs_ex_1;
input 	prifrs_ex_0;
input 	prifrs_ex_3;
input 	prifrs_ex_2;
input 	prifrs_ex_4;
output 	always02;
output 	ptAScr;
input 	always03;
output 	exmem_en;
input 	Equal1;
input 	ccifiwait_0;
output 	always1;
output 	ifid_en;
output 	pc_en;
output 	flush_idex;
input 	prifhalt_wb;
output 	ifid_en1;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \always1~1_combout ;
wire \always1~2_combout ;
wire \Equal1~0_combout ;
wire \ptBScr~0_combout ;
wire \Equal5~0_combout ;
wire \Equal4~2_combout ;
wire \Equal4~3_combout ;
wire \Equal4~5_combout ;
wire \always0~2_combout ;
wire \Equal4~4_combout ;
wire \always0~3_combout ;
wire \always0~1_combout ;
wire \always0~4_combout ;
wire \always0~0_combout ;
wire \Equal3~0_combout ;
wire \Equal2~1_combout ;
wire \Equal2~0_combout ;
wire \Equal2~2_combout ;
wire \ptAScr~1_combout ;
wire \ptAScr~0_combout ;
wire \ptAScr~2_combout ;
wire \always0~7_combout ;
wire \always0~8_combout ;
wire \ptAScr~3_combout ;
wire \always1~0_combout ;
wire \always1~3_combout ;
wire \always1~4_combout ;
wire \always1~6_combout ;


// Location: LCCOMB_X54_Y30_N30
cycloneive_lcell_comb \always1~1 (
// Equation(s):
// \always1~1_combout  = (!\prif.opcode_mem [0] & (!\prif.instr_mem [4] & (!\prif.instr_mem [5] & \prif.instr_mem [3])))

	.dataa(prifopcode_mem_0),
	.datab(prifinstr_mem_4),
	.datac(prifinstr_mem_5),
	.datad(prifinstr_mem_3),
	.cin(gnd),
	.combout(\always1~1_combout ),
	.cout());
// synopsys translate_off
defparam \always1~1 .lut_mask = 16'h0100;
defparam \always1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N20
cycloneive_lcell_comb \always1~2 (
// Equation(s):
// \always1~2_combout  = (!\prif.instr_mem [1] & (!\prif.instr_mem [2] & (\always1~1_combout  & !\prif.instr_mem [0])))

	.dataa(prifinstr_mem_1),
	.datab(prifinstr_mem_2),
	.datac(\always1~1_combout ),
	.datad(prifinstr_mem_0),
	.cin(gnd),
	.combout(\always1~2_combout ),
	.cout());
// synopsys translate_off
defparam \always1~2 .lut_mask = 16'h0010;
defparam \always1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N16
cycloneive_lcell_comb \ptBScr~1 (
// Equation(s):
// ptBScr = (\ptBScr~0_combout  & (\Equal4~5_combout  & ((\prif.rt_ex [4]) # (!\Equal5~0_combout ))))

	.dataa(\ptBScr~0_combout ),
	.datab(prifrt_ex_4),
	.datac(\Equal5~0_combout ),
	.datad(\Equal4~5_combout ),
	.cin(gnd),
	.combout(ptBScr),
	.cout());
// synopsys translate_off
defparam \ptBScr~1 .lut_mask = 16'h8A00;
defparam \ptBScr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N20
cycloneive_lcell_comb \Equal8~0 (
// Equation(s):
// Equal8 = (!\prif.regwrite_wb [3] & (!\prif.regwrite_wb [1] & !\prif.regwrite_wb [4]))

	.dataa(gnd),
	.datab(prifregwrite_wb_3),
	.datac(prifregwrite_wb_1),
	.datad(prifregwrite_wb_4),
	.cin(gnd),
	.combout(Equal8),
	.cout());
// synopsys translate_off
defparam \Equal8~0 .lut_mask = 16'h0003;
defparam \Equal8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N20
cycloneive_lcell_comb \always0~5 (
// Equation(s):
// always01 = (\always0~3_combout  & (\always0~1_combout  & (\always0~4_combout  & \always0~0_combout )))

	.dataa(\always0~3_combout ),
	.datab(\always0~1_combout ),
	.datac(\always0~4_combout ),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(always01),
	.cout());
// synopsys translate_off
defparam \always0~5 .lut_mask = 16'h8000;
defparam \always0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N0
cycloneive_lcell_comb \always0~6 (
// Equation(s):
// always02 = (\ptBScr~0_combout  & (\Equal2~2_combout  & ((\prif.rs_ex [0]) # (!\Equal3~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(prifrs_ex_0),
	.datac(\ptBScr~0_combout ),
	.datad(\Equal2~2_combout ),
	.cin(gnd),
	.combout(always02),
	.cout());
// synopsys translate_off
defparam \always0~6 .lut_mask = 16'hD000;
defparam \always0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N14
cycloneive_lcell_comb \ptAScr~4 (
// Equation(s):
// ptAScr = (\ptAScr~2_combout  & (always02 & (\always0~8_combout ))) # (!\ptAScr~2_combout  & (((\ptAScr~3_combout ))))

	.dataa(\ptAScr~2_combout ),
	.datab(always02),
	.datac(\always0~8_combout ),
	.datad(\ptAScr~3_combout ),
	.cin(gnd),
	.combout(ptAScr),
	.cout());
// synopsys translate_off
defparam \ptAScr~4 .lut_mask = 16'hD580;
defparam \ptAScr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N26
cycloneive_lcell_comb \exmem_en~0 (
// Equation(s):
// exmem_en = (!always01 & (((LessThan1 & always0)) # (!\nRST~input_o )))

	.dataa(nRST),
	.datab(LessThan1),
	.datac(always0),
	.datad(always03),
	.cin(gnd),
	.combout(exmem_en),
	.cout());
// synopsys translate_off
defparam \exmem_en~0 .lut_mask = 16'h00D5;
defparam \exmem_en~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N22
cycloneive_lcell_comb \always1~5 (
// Equation(s):
// always1 = (!ccifiwait_0 & ((\always1~4_combout ) # ((\Equal1~1_combout  & \prif.zero_flag_mem~q ))))

	.dataa(Equal1),
	.datab(ccifiwait_0),
	.datac(prifzero_flag_mem),
	.datad(\always1~4_combout ),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~5 .lut_mask = 16'h3320;
defparam \always1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N14
cycloneive_lcell_comb \ifid_en~0 (
// Equation(s):
// ifid_en = (((ccifiwait_0) # (always1)) # (!\prif.opcode_ex [5])) # (!\always1~6_combout )

	.dataa(\always1~6_combout ),
	.datab(prifopcode_ex_5),
	.datac(ccifiwait_0),
	.datad(always1),
	.cin(gnd),
	.combout(ifid_en),
	.cout());
// synopsys translate_off
defparam \ifid_en~0 .lut_mask = 16'hFFF7;
defparam \ifid_en~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N6
cycloneive_lcell_comb \pc_en~0 (
// Equation(s):
// pc_en = (exmem_en & ifid_en)

	.dataa(exmem_en),
	.datab(gnd),
	.datac(ifid_en),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_en),
	.cout());
// synopsys translate_off
defparam \pc_en~0 .lut_mask = 16'hA0A0;
defparam \pc_en~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N24
cycloneive_lcell_comb \flush_idex~0 (
// Equation(s):
// flush_idex = (always1) # ((\always1~6_combout  & (!ccifiwait_0 & \prif.opcode_ex [5])))

	.dataa(\always1~6_combout ),
	.datab(ccifiwait_0),
	.datac(prifopcode_ex_5),
	.datad(always1),
	.cin(gnd),
	.combout(flush_idex),
	.cout());
// synopsys translate_off
defparam \flush_idex~0 .lut_mask = 16'hFF20;
defparam \flush_idex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N10
cycloneive_lcell_comb \ifid_en~1 (
// Equation(s):
// ifid_en1 = (!ccifiwait_0 & (ifid_en & !\prif.halt_wb~q ))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(ifid_en),
	.datad(prifhalt_wb),
	.cin(gnd),
	.combout(ifid_en1),
	.cout());
// synopsys translate_off
defparam \ifid_en~1 .lut_mask = 16'h0030;
defparam \ifid_en~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N8
cycloneive_lcell_comb \Equal1~0 (
// Equation(s):
// \Equal1~0_combout  = (!\prif.regwrite_mem [3] & (!\prif.regwrite_mem [0] & (!\prif.regwrite_mem [1] & !\prif.regwrite_mem [2])))

	.dataa(prifregwrite_mem_3),
	.datab(prifregwrite_mem_0),
	.datac(prifregwrite_mem_1),
	.datad(prifregwrite_mem_2),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0001;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N30
cycloneive_lcell_comb \ptBScr~0 (
// Equation(s):
// \ptBScr~0_combout  = (\prif.Regwen_mem~q  & ((\prif.regwrite_mem [4]) # (!\Equal1~0_combout )))

	.dataa(prifRegwen_mem),
	.datab(gnd),
	.datac(\Equal1~0_combout ),
	.datad(prifregwrite_mem_4),
	.cin(gnd),
	.combout(\ptBScr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ptBScr~0 .lut_mask = 16'hAA0A;
defparam \ptBScr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N22
cycloneive_lcell_comb \Equal5~0 (
// Equation(s):
// \Equal5~0_combout  = (!\prif.rt_ex [2] & (!\prif.rt_ex [1] & (!\prif.rt_ex [3] & !\prif.rt_ex [0])))

	.dataa(prifrt_ex_2),
	.datab(prifrt_ex_1),
	.datac(prifrt_ex_3),
	.datad(prifrt_ex_0),
	.cin(gnd),
	.combout(\Equal5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal5~0 .lut_mask = 16'h0001;
defparam \Equal5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N26
cycloneive_lcell_comb \Equal4~2 (
// Equation(s):
// \Equal4~2_combout  = (\prif.regwrite_mem [0] & (\prif.rt_ex [0] & (\prif.rt_ex [1] $ (!\prif.regwrite_mem [1])))) # (!\prif.regwrite_mem [0] & (!\prif.rt_ex [0] & (\prif.rt_ex [1] $ (!\prif.regwrite_mem [1]))))

	.dataa(prifregwrite_mem_0),
	.datab(prifrt_ex_0),
	.datac(prifrt_ex_1),
	.datad(prifregwrite_mem_1),
	.cin(gnd),
	.combout(\Equal4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~2 .lut_mask = 16'h9009;
defparam \Equal4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N0
cycloneive_lcell_comb \Equal4~3 (
// Equation(s):
// \Equal4~3_combout  = (\prif.rt_ex [2] & (\prif.regwrite_mem [2] & (\prif.rt_ex [3] $ (!\prif.regwrite_mem [3])))) # (!\prif.rt_ex [2] & (!\prif.regwrite_mem [2] & (\prif.rt_ex [3] $ (!\prif.regwrite_mem [3]))))

	.dataa(prifrt_ex_2),
	.datab(prifrt_ex_3),
	.datac(prifregwrite_mem_2),
	.datad(prifregwrite_mem_3),
	.cin(gnd),
	.combout(\Equal4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~3 .lut_mask = 16'h8421;
defparam \Equal4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N18
cycloneive_lcell_comb \Equal4~5 (
// Equation(s):
// \Equal4~5_combout  = (\Equal4~2_combout  & (\Equal4~3_combout  & (\prif.rt_ex [4] $ (!\prif.regwrite_mem [4]))))

	.dataa(\Equal4~2_combout ),
	.datab(prifrt_ex_4),
	.datac(prifregwrite_mem_4),
	.datad(\Equal4~3_combout ),
	.cin(gnd),
	.combout(\Equal4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~5 .lut_mask = 16'h8200;
defparam \Equal4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N30
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// \always0~2_combout  = (\prif.rt_ex [2] & (\prif.regwrite_wb [2] & (\prif.regwrite_wb [3] $ (!\prif.rt_ex [3])))) # (!\prif.rt_ex [2] & (!\prif.regwrite_wb [2] & (\prif.regwrite_wb [3] $ (!\prif.rt_ex [3]))))

	.dataa(prifrt_ex_2),
	.datab(prifregwrite_wb_3),
	.datac(prifrt_ex_3),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'h8241;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N16
cycloneive_lcell_comb \Equal4~4 (
// Equation(s):
// \Equal4~4_combout  = \prif.rt_ex [4] $ (\prif.regwrite_mem [4])

	.dataa(prifrt_ex_4),
	.datab(gnd),
	.datac(gnd),
	.datad(prifregwrite_mem_4),
	.cin(gnd),
	.combout(\Equal4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Equal4~4 .lut_mask = 16'h55AA;
defparam \Equal4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N12
cycloneive_lcell_comb \always0~3 (
// Equation(s):
// \always0~3_combout  = (\always0~2_combout  & (((\Equal4~4_combout ) # (!\Equal4~3_combout )) # (!\Equal4~2_combout )))

	.dataa(\Equal4~2_combout ),
	.datab(\Equal4~3_combout ),
	.datac(\always0~2_combout ),
	.datad(\Equal4~4_combout ),
	.cin(gnd),
	.combout(\always0~3_combout ),
	.cout());
// synopsys translate_off
defparam \always0~3 .lut_mask = 16'hF070;
defparam \always0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N28
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (\prif.rt_ex [1] & (\prif.regwrite_wb [1] & (\prif.regwrite_wb [0] $ (!\prif.rt_ex [0])))) # (!\prif.rt_ex [1] & (!\prif.regwrite_wb [1] & (\prif.regwrite_wb [0] $ (!\prif.rt_ex [0]))))

	.dataa(prifrt_ex_1),
	.datab(prifregwrite_wb_0),
	.datac(prifregwrite_wb_1),
	.datad(prifrt_ex_0),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'h8421;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N14
cycloneive_lcell_comb \always0~4 (
// Equation(s):
// \always0~4_combout  = (\prif.regwrite_wb [4] & (\prif.rt_ex [4])) # (!\prif.regwrite_wb [4] & (!\prif.rt_ex [4] & !\Equal5~0_combout ))

	.dataa(prifregwrite_wb_4),
	.datab(prifrt_ex_4),
	.datac(\Equal5~0_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\always0~4_combout ),
	.cout());
// synopsys translate_off
defparam \always0~4 .lut_mask = 16'h8989;
defparam \always0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N6
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (\prif.Regwen_wb~q  & ((\prif.regwrite_wb [0]) # ((\prif.regwrite_wb [2]) # (!Equal8))))

	.dataa(prifRegwen_wb),
	.datab(prifregwrite_wb_0),
	.datac(Equal8),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'hAA8A;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N10
cycloneive_lcell_comb \Equal3~0 (
// Equation(s):
// \Equal3~0_combout  = (!\prif.rs_ex [1] & (!\prif.rs_ex [3] & (!\prif.rs_ex [2] & !\prif.rs_ex [4])))

	.dataa(prifrs_ex_1),
	.datab(prifrs_ex_3),
	.datac(prifrs_ex_2),
	.datad(prifrs_ex_4),
	.cin(gnd),
	.combout(\Equal3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal3~0 .lut_mask = 16'h0001;
defparam \Equal3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N8
cycloneive_lcell_comb \Equal2~1 (
// Equation(s):
// \Equal2~1_combout  = (\prif.regwrite_mem [3] & (\prif.rs_ex [3] & (\prif.regwrite_mem [2] $ (!\prif.rs_ex [2])))) # (!\prif.regwrite_mem [3] & (!\prif.rs_ex [3] & (\prif.regwrite_mem [2] $ (!\prif.rs_ex [2]))))

	.dataa(prifregwrite_mem_3),
	.datab(prifregwrite_mem_2),
	.datac(prifrs_ex_2),
	.datad(prifrs_ex_3),
	.cin(gnd),
	.combout(\Equal2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~1 .lut_mask = 16'h8241;
defparam \Equal2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N2
cycloneive_lcell_comb \Equal2~0 (
// Equation(s):
// \Equal2~0_combout  = (\prif.rs_ex [1] & (\prif.regwrite_mem [1] & (\prif.rs_ex [0] $ (!\prif.regwrite_mem [0])))) # (!\prif.rs_ex [1] & (!\prif.regwrite_mem [1] & (\prif.rs_ex [0] $ (!\prif.regwrite_mem [0]))))

	.dataa(prifrs_ex_1),
	.datab(prifrs_ex_0),
	.datac(prifregwrite_mem_1),
	.datad(prifregwrite_mem_0),
	.cin(gnd),
	.combout(\Equal2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~0 .lut_mask = 16'h8421;
defparam \Equal2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N24
cycloneive_lcell_comb \Equal2~2 (
// Equation(s):
// \Equal2~2_combout  = (\Equal2~1_combout  & (\Equal2~0_combout  & (\prif.rs_ex [4] $ (!\prif.regwrite_mem [4]))))

	.dataa(prifrs_ex_4),
	.datab(prifregwrite_mem_4),
	.datac(\Equal2~1_combout ),
	.datad(\Equal2~0_combout ),
	.cin(gnd),
	.combout(\Equal2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Equal2~2 .lut_mask = 16'h9000;
defparam \Equal2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N4
cycloneive_lcell_comb \ptAScr~1 (
// Equation(s):
// \ptAScr~1_combout  = (\prif.rs_ex [4] & ((\prif.regwrite_wb [1] $ (\prif.rs_ex [1])) # (!\prif.regwrite_wb [4]))) # (!\prif.rs_ex [4] & ((\prif.regwrite_wb [4]) # (\prif.regwrite_wb [1] $ (\prif.rs_ex [1]))))

	.dataa(prifrs_ex_4),
	.datab(prifregwrite_wb_1),
	.datac(prifrs_ex_1),
	.datad(prifregwrite_wb_4),
	.cin(gnd),
	.combout(\ptAScr~1_combout ),
	.cout());
// synopsys translate_off
defparam \ptAScr~1 .lut_mask = 16'h7DBE;
defparam \ptAScr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N18
cycloneive_lcell_comb \ptAScr~0 (
// Equation(s):
// \ptAScr~0_combout  = (\prif.regwrite_wb [3] & ((\prif.regwrite_wb [2] $ (\prif.rs_ex [2])) # (!\prif.rs_ex [3]))) # (!\prif.regwrite_wb [3] & ((\prif.rs_ex [3]) # (\prif.regwrite_wb [2] $ (\prif.rs_ex [2]))))

	.dataa(prifregwrite_wb_3),
	.datab(prifregwrite_wb_2),
	.datac(prifrs_ex_2),
	.datad(prifrs_ex_3),
	.cin(gnd),
	.combout(\ptAScr~0_combout ),
	.cout());
// synopsys translate_off
defparam \ptAScr~0 .lut_mask = 16'h7DBE;
defparam \ptAScr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N22
cycloneive_lcell_comb \ptAScr~2 (
// Equation(s):
// \ptAScr~2_combout  = (\ptAScr~1_combout ) # ((\ptAScr~0_combout ) # (\prif.regwrite_wb [0] $ (\prif.rs_ex [0])))

	.dataa(prifregwrite_wb_0),
	.datab(prifrs_ex_0),
	.datac(\ptAScr~1_combout ),
	.datad(\ptAScr~0_combout ),
	.cin(gnd),
	.combout(\ptAScr~2_combout ),
	.cout());
// synopsys translate_off
defparam \ptAScr~2 .lut_mask = 16'hFFF6;
defparam \ptAScr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N22
cycloneive_lcell_comb \always0~7 (
// Equation(s):
// \always0~7_combout  = (\prif.opcode_mem [2] & (!\prif.opcode_mem [5] & (!\prif.opcode_mem [4] & \prif.opcode_mem [3])))

	.dataa(prifopcode_mem_2),
	.datab(prifopcode_mem_5),
	.datac(prifopcode_mem_4),
	.datad(prifopcode_mem_3),
	.cin(gnd),
	.combout(\always0~7_combout ),
	.cout());
// synopsys translate_off
defparam \always0~7 .lut_mask = 16'h0200;
defparam \always0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N4
cycloneive_lcell_comb \always0~8 (
// Equation(s):
// \always0~8_combout  = (\prif.opcode_mem [1] & (\always0~7_combout  & \prif.opcode_mem [0]))

	.dataa(gnd),
	.datab(prifopcode_mem_1),
	.datac(\always0~7_combout ),
	.datad(prifopcode_mem_0),
	.cin(gnd),
	.combout(\always0~8_combout ),
	.cout());
// synopsys translate_off
defparam \always0~8 .lut_mask = 16'hC000;
defparam \always0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N12
cycloneive_lcell_comb \ptAScr~3 (
// Equation(s):
// \ptAScr~3_combout  = (!\Equal2~2_combout  & (\always0~0_combout  & ((\prif.regwrite_wb [0]) # (!\Equal3~0_combout ))))

	.dataa(\Equal3~0_combout ),
	.datab(\Equal2~2_combout ),
	.datac(prifregwrite_wb_0),
	.datad(\always0~0_combout ),
	.cin(gnd),
	.combout(\ptAScr~3_combout ),
	.cout());
// synopsys translate_off
defparam \ptAScr~3 .lut_mask = 16'h3100;
defparam \ptAScr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N0
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// \always1~0_combout  = (!\prif.zero_flag_mem~q  & (!\prif.opcode_mem [1] & (\prif.opcode_mem [2] & \prif.opcode_mem [0])))

	.dataa(prifzero_flag_mem),
	.datab(prifopcode_mem_1),
	.datac(prifopcode_mem_2),
	.datad(prifopcode_mem_0),
	.cin(gnd),
	.combout(\always1~0_combout ),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'h1000;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N26
cycloneive_lcell_comb \always1~3 (
// Equation(s):
// \always1~3_combout  = (\always1~0_combout ) # ((!\prif.opcode_mem [2] & ((\always1~2_combout ) # (\prif.opcode_mem [1]))))

	.dataa(\always1~2_combout ),
	.datab(prifopcode_mem_1),
	.datac(prifopcode_mem_2),
	.datad(\always1~0_combout ),
	.cin(gnd),
	.combout(\always1~3_combout ),
	.cout());
// synopsys translate_off
defparam \always1~3 .lut_mask = 16'hFF0E;
defparam \always1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N18
cycloneive_lcell_comb \always1~4 (
// Equation(s):
// \always1~4_combout  = (!\prif.opcode_mem [4] & (!\prif.opcode_mem [5] & (\always1~3_combout  & !\prif.opcode_mem [3])))

	.dataa(prifopcode_mem_4),
	.datab(prifopcode_mem_5),
	.datac(\always1~3_combout ),
	.datad(prifopcode_mem_3),
	.cin(gnd),
	.combout(\always1~4_combout ),
	.cout());
// synopsys translate_off
defparam \always1~4 .lut_mask = 16'h0010;
defparam \always1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N14
cycloneive_lcell_comb \always1~6 (
// Equation(s):
// \always1~6_combout  = (!\prif.opcode_ex [2] & (\prif.opcode_ex [0] & (\prif.opcode_ex [1] & !\prif.opcode_ex [4])))

	.dataa(prifopcode_ex_2),
	.datab(prifopcode_ex_0),
	.datac(prifopcode_ex_1),
	.datad(prifopcode_ex_4),
	.cin(gnd),
	.combout(\always1~6_combout ),
	.cout());
// synopsys translate_off
defparam \always1~6 .lut_mask = 16'h0040;
defparam \always1~6 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module pipeline_register (
	prifdmemaddr_1,
	pc_1,
	prifdmemren,
	prifdmemwen,
	prifdmemaddr_0,
	pc_0,
	prifdmemaddr_3,
	prifdmemaddr_2,
	prifdmemaddr_5,
	prifdmemaddr_4,
	prifdmemaddr_7,
	prifdmemaddr_6,
	prifdmemaddr_9,
	prifdmemaddr_8,
	prifdmemaddr_11,
	prifdmemaddr_10,
	prifdmemaddr_13,
	prifdmemaddr_12,
	prifdmemaddr_15,
	prifdmemaddr_14,
	prifdmemaddr_23,
	prifdmemaddr_22,
	prifdmemaddr_21,
	prifdmemaddr_29,
	prifdmemaddr_28,
	prifdmemaddr_31,
	prifdmemaddr_30,
	prifdmemaddr_20,
	prifdmemaddr_17,
	prifdmemaddr_16,
	prifdmemaddr_19,
	prifdmemaddr_18,
	prifdmemaddr_25,
	prifdmemaddr_24,
	prifdmemaddr_27,
	prifdmemaddr_26,
	prifhalt_mem,
	prifdmemstore_0,
	prifimm_ex_1,
	prifALUScr_ex_1,
	prifshamt_ex_1,
	prifALUScr_ex_0,
	prifRegwen_mem,
	prifregwrite_mem_4,
	prifregwrite_mem_0,
	prifregwrite_mem_1,
	prifregwrite_mem_2,
	prifregwrite_mem_3,
	prifrt_ex_1,
	prifrt_ex_0,
	prifrt_ex_3,
	prifrt_ex_2,
	prifrt_ex_4,
	prifrdat2_ex_1,
	prifopcode_mem_1,
	prifopcode_mem_0,
	prifopcode_mem_2,
	prifopcode_mem_3,
	prifopcode_mem_5,
	prifopcode_mem_4,
	prifrdat1_ex_1,
	prifimm_ex_0,
	prifshamt_ex_0,
	prifrdat2_ex_0,
	prifrdat1_ex_0,
	prifrdat2_ex_3,
	prifimm_ex_3,
	prifshamt_ex_3,
	prifimm_ex_2,
	prifshamt_ex_2,
	prifrdat2_ex_2,
	prifrdat2_ex_4,
	prifimm_ex_4,
	prifshamt_ex_4,
	prifinstr_ex_15,
	prifrdat2_ex_31,
	prifimm_mem_15,
	prifrdat2_ex_30,
	prifimm_mem_14,
	prifrdat2_ex_29,
	prifimm_mem_13,
	prifimm_ex_5,
	prifrdat2_ex_5,
	prifimm_ex_15,
	prifrdat2_ex_15,
	prifimm_ex_14,
	prifrdat2_ex_14,
	prifimm_ex_13,
	prifrdat2_ex_13,
	prifimm_ex_12,
	prifrdat2_ex_12,
	prifimm_ex_11,
	prifrdat2_ex_11,
	prifimm_ex_10,
	prifrdat2_ex_10,
	prifimm_ex_9,
	prifrdat2_ex_9,
	prifimm_ex_6,
	prifrdat2_ex_6,
	prifrdat2_ex_27,
	prifimm_mem_11,
	prifrdat2_ex_23,
	prifimm_mem_7,
	prifrdat2_ex_18,
	prifimm_mem_2,
	prifrdat2_ex_24,
	prifimm_mem_8,
	prifrdat2_ex_16,
	prifimm_mem_0,
	prifrdat2_ex_19,
	prifimm_mem_3,
	prifrdat2_ex_17,
	prifimm_mem_1,
	prifrdat2_ex_21,
	prifimm_mem_5,
	prifrdat2_ex_20,
	prifimm_mem_4,
	prifrdat2_ex_28,
	prifimm_mem_12,
	prifrdat2_ex_26,
	prifimm_mem_10,
	prifimm_ex_8,
	prifrdat2_ex_8,
	prifimm_ex_7,
	prifrdat2_ex_7,
	prifrdat2_ex_22,
	prifimm_mem_6,
	prifrdat2_ex_25,
	prifimm_mem_9,
	prifrdat1_ex_2,
	prifrdat1_ex_4,
	prifrdat1_ex_3,
	prifrdat1_ex_8,
	prifrdat1_ex_7,
	prifrdat1_ex_6,
	prifrdat1_ex_5,
	prifrdat1_ex_16,
	prifrdat1_ex_15,
	prifrdat1_ex_14,
	prifrdat1_ex_13,
	prifrdat1_ex_11,
	prifrdat1_ex_12,
	prifrdat1_ex_10,
	prifrdat1_ex_9,
	prifrdat1_ex_18,
	prifrdat1_ex_17,
	prifrdat1_ex_20,
	prifrdat1_ex_19,
	prifrdat1_ex_22,
	prifrdat1_ex_21,
	prifrdat1_ex_24,
	prifrdat1_ex_23,
	prifrdat1_ex_31,
	prifrdat1_ex_30,
	prifrdat1_ex_29,
	prifrdat1_ex_26,
	prifrdat1_ex_25,
	prifrdat1_ex_28,
	prifrdat1_ex_27,
	prifzero_flag_mem,
	prifinstr_mem_3,
	prifinstr_mem_5,
	prifinstr_mem_4,
	prifinstr_mem_2,
	prifinstr_mem_1,
	prifinstr_mem_0,
	prifrdat1_mem_1,
	prifPCScr_mem_0,
	prifpc_bran_mem_1,
	prifPCScr_mem_1,
	prifopcode_ex_5,
	prifopcode_ex_0,
	prifopcode_ex_1,
	prifopcode_ex_2,
	prifopcode_ex_4,
	prifmemren_ex,
	prifmemwen_ex,
	prifrdat1_mem_0,
	prifpc_bran_mem_0,
	prifrdat1_mem_3,
	prifpc_bran_mem_3,
	prifrdat1_mem_2,
	prifpc_bran_mem_2,
	prifrdat1_mem_5,
	prifpc_bran_mem_5,
	prifrdat1_mem_4,
	prifpc_bran_mem_4,
	prifrdat1_mem_7,
	prifpc_bran_mem_7,
	prifrdat1_mem_6,
	prifpc_bran_mem_6,
	prifrdat1_mem_9,
	prifpc_bran_mem_9,
	prifinstr_mem_7,
	prifrdat1_mem_8,
	prifpc_bran_mem_8,
	prifinstr_mem_6,
	prifrdat1_mem_11,
	prifpc_bran_mem_11,
	prifinstr_mem_9,
	prifrdat1_mem_10,
	prifpc_bran_mem_10,
	prifinstr_mem_8,
	prifrdat1_mem_13,
	prifpc_bran_mem_13,
	prifinstr_mem_11,
	prifrdat1_mem_12,
	prifpc_bran_mem_12,
	prifinstr_mem_10,
	prifrdat1_mem_15,
	prifpc_bran_mem_15,
	prifinstr_mem_13,
	prifrdat1_mem_14,
	prifpc_bran_mem_14,
	prifinstr_mem_12,
	prifrdat1_mem_23,
	prifpc_bran_mem_23,
	prifinstr_mem_21,
	prifrdat1_mem_22,
	prifpc_bran_mem_22,
	prifinstr_mem_20,
	prifrdat1_mem_21,
	prifpc_bran_mem_21,
	prifinstr_mem_19,
	prifrdat1_mem_29,
	prifpc_bran_mem_29,
	prifrdat1_mem_28,
	prifpc_bran_mem_28,
	prifrdat1_mem_31,
	prifpc_bran_mem_31,
	prifrdat1_mem_30,
	prifpc_bran_mem_30,
	prifrdat1_mem_20,
	prifpc_bran_mem_20,
	prifinstr_mem_18,
	prifrdat1_mem_17,
	prifpc_bran_mem_17,
	prifinstr_mem_15,
	prifrdat1_mem_16,
	prifpc_bran_mem_16,
	prifinstr_mem_14,
	prifrdat1_mem_19,
	prifpc_bran_mem_19,
	prifinstr_mem_17,
	prifrdat1_mem_18,
	prifpc_bran_mem_18,
	prifinstr_mem_16,
	prifrdat1_mem_25,
	prifpc_bran_mem_25,
	prifinstr_mem_23,
	prifrdat1_mem_24,
	prifpc_bran_mem_24,
	prifinstr_mem_22,
	prifrdat1_mem_27,
	prifpc_bran_mem_27,
	prifinstr_mem_25,
	prifrdat1_mem_26,
	prifpc_bran_mem_26,
	prifinstr_mem_24,
	prifdmemstore_1,
	prifdmemstore_2,
	prifdmemstore_3,
	prifdmemstore_4,
	prifdmemstore_5,
	prifdmemstore_6,
	prifdmemstore_7,
	prifdmemstore_8,
	prifdmemstore_9,
	prifdmemstore_10,
	prifdmemstore_11,
	prifdmemstore_12,
	prifdmemstore_13,
	prifdmemstore_14,
	prifdmemstore_15,
	prifdmemstore_16,
	prifdmemstore_17,
	prifdmemstore_18,
	prifdmemstore_19,
	prifdmemstore_20,
	prifdmemstore_21,
	prifdmemstore_22,
	prifdmemstore_23,
	prifdmemstore_24,
	prifdmemstore_25,
	prifdmemstore_26,
	prifdmemstore_27,
	prifdmemstore_28,
	prifdmemstore_29,
	prifdmemstore_30,
	prifdmemstore_31,
	prifhalt_ex,
	prifimemload_id_31,
	prifimemload_id_30,
	prifimemload_id_29,
	prifimemload_id_27,
	prifimemload_id_26,
	prifimemload_id_28,
	prifimemload_id_3,
	prifimemload_id_1,
	prifimemload_id_5,
	prifimemload_id_4,
	prifimemload_id_2,
	prifimemload_id_0,
	prifimemload_id_7,
	prifRegwen_ex,
	prifrd_ex_4,
	prifRegDest_ex_1,
	prifRegDest_ex_0,
	prifrd_ex_0,
	prifrd_ex_1,
	prifrd_ex_2,
	prifrd_ex_3,
	prifimemload_id_17,
	prifimemload_id_16,
	prifimemload_id_19,
	prifimemload_id_18,
	prifimemload_id_20,
	prifdataScr_mem_0,
	prifdataScr_mem_1,
	prifimemload_id_22,
	prifimemload_id_21,
	prifimemload_id_24,
	prifimemload_id_23,
	prifimemload_id_25,
	prifopcode_ex_3,
	prifimemload_id_6,
	prifimemload_id_9,
	prifimemload_id_8,
	prifimemload_id_10,
	prifimemload_id_15,
	prifimemload_id_14,
	prifimemload_id_13,
	prifimemload_id_12,
	prifimemload_id_11,
	prifinstr_ex_3,
	prifinstr_ex_5,
	prifinstr_ex_4,
	prifinstr_ex_2,
	prifinstr_ex_1,
	prifinstr_ex_0,
	prifPCScr_ex_0,
	prifpc_ex_1,
	prifPCScr_ex_1,
	prifpc_ex_0,
	prifpc_ex_3,
	prifpc_ex_2,
	Add0,
	Add01,
	prifpc_ex_5,
	prifpc_ex_4,
	Add02,
	Add03,
	prifpc_ex_7,
	prifpc_ex_6,
	Add04,
	Add05,
	prifpc_ex_9,
	prifpc_ex_8,
	Add06,
	Add07,
	prifinstr_ex_7,
	prifinstr_ex_6,
	prifpc_ex_11,
	prifpc_ex_10,
	Add08,
	Add09,
	prifinstr_ex_9,
	prifinstr_ex_8,
	prifpc_ex_13,
	prifpc_ex_12,
	Add010,
	Add011,
	prifinstr_ex_11,
	prifinstr_ex_10,
	prifpc_ex_15,
	prifpc_ex_14,
	Add012,
	Add013,
	prifinstr_ex_13,
	prifinstr_ex_12,
	prifpc_ex_23,
	prifpc_ex_22,
	prifpc_ex_21,
	prifpc_ex_20,
	prifpc_ex_19,
	prifpc_ex_18,
	prifpc_ex_17,
	prifpc_ex_16,
	Add014,
	Add015,
	Add016,
	Add017,
	Add018,
	Add019,
	Add020,
	Add021,
	prifinstr_ex_21,
	prifinstr_ex_20,
	prifinstr_ex_19,
	prifpc_ex_29,
	prifpc_ex_28,
	prifpc_ex_27,
	prifpc_ex_26,
	prifpc_ex_25,
	prifpc_ex_24,
	Add022,
	Add023,
	Add024,
	Add025,
	Add026,
	Add027,
	prifpc_ex_31,
	prifpc_ex_30,
	Add028,
	Add029,
	prifinstr_ex_18,
	prifinstr_ex_14,
	prifinstr_ex_17,
	prifinstr_ex_16,
	prifinstr_ex_23,
	prifinstr_ex_22,
	prifinstr_ex_25,
	prifinstr_ex_24,
	prifdataScr_ex_0,
	prifdataScr_ex_1,
	prifpc_id_1,
	prifpc_id_0,
	prifpc_id_3,
	prifpc_id_2,
	prifpc_id_5,
	prifpc_id_4,
	prifpc_id_7,
	prifpc_id_6,
	prifpc_id_9,
	prifpc_id_8,
	prifpc_id_11,
	prifpc_id_10,
	prifpc_id_13,
	prifpc_id_12,
	prifpc_id_15,
	prifpc_id_14,
	prifpc_id_23,
	prifpc_id_22,
	prifpc_id_21,
	prifpc_id_20,
	prifpc_id_19,
	prifpc_id_18,
	prifpc_id_17,
	prifpc_id_16,
	prifpc_id_29,
	prifpc_id_28,
	prifpc_id_27,
	prifpc_id_26,
	prifpc_id_25,
	prifpc_id_24,
	prifpc_id_31,
	prifpc_id_30,
	Add2,
	Add21,
	Add22,
	Add23,
	Add24,
	Add25,
	Add26,
	Add27,
	Add28,
	Add29,
	Add210,
	Add211,
	Add212,
	Add213,
	Add214,
	Add215,
	Add216,
	Add217,
	Add218,
	Add219,
	Add220,
	Add221,
	Add222,
	Add223,
	Add224,
	Add225,
	Add226,
	Add227,
	Add228,
	pc_2,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	prifALUOP_ex_3,
	prifRegwen_wb,
	prifregwrite_wb_2,
	prifregwrite_wb_0,
	prifregwrite_wb_1,
	prifregwrite_wb_4,
	prifregwrite_wb_3,
	Mux62,
	prifdmemload_wb_1,
	prifdmemaddr_wb_1,
	prifdataScr_wb_0,
	prifdataScr_wb_1,
	prifpc_wb_1,
	Mux621,
	prifrs_ex_1,
	prifrs_ex_0,
	prifrs_ex_3,
	prifrs_ex_2,
	prifrs_ex_4,
	Mux63,
	prifdmemload_wb_0,
	prifdmemaddr_wb_0,
	prifpc_wb_0,
	Mux631,
	prifdmemload_wb_3,
	prifdmemaddr_wb_3,
	prifpc_wb_3,
	prifdmemload_wb_2,
	prifdmemaddr_wb_2,
	prifpc_wb_2,
	Mux61,
	prifdmemload_wb_4,
	prifdmemaddr_wb_4,
	prifpc_wb_4,
	prifdmemload_wb_31,
	prifimm_wb_15,
	prifdmemaddr_wb_31,
	prifpc_wb_31,
	Mux32,
	prifimm_wb_14,
	prifdmemload_wb_30,
	prifdmemaddr_wb_30,
	prifpc_wb_30,
	Mux33,
	prifdmemload_wb_29,
	prifimm_wb_13,
	prifdmemaddr_wb_29,
	prifpc_wb_29,
	Mux34,
	prifdmemload_wb_5,
	prifdmemaddr_wb_5,
	prifpc_wb_5,
	prifdmemload_wb_15,
	prifdmemaddr_wb_15,
	prifpc_wb_15,
	prifdmemload_wb_14,
	prifdmemaddr_wb_14,
	prifpc_wb_14,
	prifdmemload_wb_13,
	prifdmemaddr_wb_13,
	prifpc_wb_13,
	prifdmemload_wb_12,
	prifdmemaddr_wb_12,
	prifpc_wb_12,
	prifdmemload_wb_11,
	prifdmemaddr_wb_11,
	prifpc_wb_11,
	prifdmemload_wb_10,
	prifdmemaddr_wb_10,
	prifpc_wb_10,
	prifdmemload_wb_9,
	prifdmemaddr_wb_9,
	prifpc_wb_9,
	prifdmemload_wb_6,
	prifdmemaddr_wb_6,
	prifpc_wb_6,
	prifdmemload_wb_27,
	prifimm_wb_11,
	prifdmemaddr_wb_27,
	prifpc_wb_27,
	Mux36,
	prifdmemload_wb_23,
	prifimm_wb_7,
	prifdmemaddr_wb_23,
	prifpc_wb_23,
	Mux40,
	prifimm_wb_2,
	prifdmemload_wb_18,
	prifdmemaddr_wb_18,
	prifpc_wb_18,
	Mux45,
	prifimm_wb_8,
	prifdmemload_wb_24,
	prifdmemaddr_wb_24,
	prifpc_wb_24,
	Mux39,
	prifimm_wb_0,
	prifdmemload_wb_16,
	prifdmemaddr_wb_16,
	prifpc_wb_16,
	Mux47,
	prifdmemload_wb_19,
	prifimm_wb_3,
	prifdmemaddr_wb_19,
	prifpc_wb_19,
	Mux44,
	prifdmemload_wb_17,
	prifimm_wb_1,
	prifdmemaddr_wb_17,
	prifpc_wb_17,
	Mux46,
	prifdmemload_wb_21,
	prifimm_wb_5,
	prifdmemaddr_wb_21,
	prifpc_wb_21,
	Mux42,
	prifimm_wb_4,
	prifdmemload_wb_20,
	prifdmemaddr_wb_20,
	prifpc_wb_20,
	Mux43,
	prifimm_wb_12,
	prifdmemload_wb_28,
	prifdmemaddr_wb_28,
	prifpc_wb_28,
	Mux35,
	prifimm_wb_10,
	prifdmemload_wb_26,
	prifdmemaddr_wb_26,
	prifpc_wb_26,
	Mux37,
	prifdmemload_wb_8,
	prifdmemaddr_wb_8,
	prifpc_wb_8,
	prifdmemload_wb_7,
	prifdmemaddr_wb_7,
	prifpc_wb_7,
	prifimm_wb_6,
	prifdmemload_wb_22,
	prifdmemaddr_wb_22,
	prifpc_wb_22,
	Mux41,
	prifdmemload_wb_25,
	prifimm_wb_9,
	prifdmemaddr_wb_25,
	prifpc_wb_25,
	Mux38,
	prifALUOP_ex_2,
	prifALUOP_ex_1,
	prifALUOP_ex_0,
	aluifportOut_1,
	exmem_en,
	dmemaddr,
	ccifiwait_0,
	dmemren,
	dmemwen,
	aluifportOut_0,
	dmemaddr1,
	aluifportOut_3,
	aluifportOut_5,
	aluifportOut_2,
	aluifportOut_31,
	aluifportOut_32,
	dmemaddr2,
	aluifportOut_21,
	dmemaddr3,
	aluifportOut_51,
	aluifportOut_52,
	dmemaddr4,
	aluifportOut_4,
	dmemaddr5,
	aluifportOut_7,
	dmemaddr6,
	aluifportOut_6,
	dmemaddr7,
	aluifportOut_9,
	dmemaddr8,
	aluifportOut_8,
	dmemaddr9,
	aluifportOut_11,
	dmemaddr10,
	aluifportOut_10,
	dmemaddr11,
	aluifportOut_13,
	dmemaddr12,
	aluifportOut_12,
	dmemaddr13,
	aluifportOut_15,
	dmemaddr14,
	aluifportOut_14,
	dmemaddr15,
	aluifportOut_23,
	dmemaddr16,
	aluifportOut_22,
	dmemaddr17,
	aluifportOut_211,
	dmemaddr18,
	aluifportOut_29,
	dmemaddr19,
	prifpc_mem_29,
	aluifportOut_28,
	dmemaddr20,
	prifpc_mem_28,
	aluifneg_flag,
	dmemaddr21,
	prifpc_mem_31,
	aluifportOut_30,
	dmemaddr22,
	prifpc_mem_30,
	aluifportOut_20,
	dmemaddr23,
	aluifportOut_17,
	dmemaddr24,
	aluifportOut_16,
	dmemaddr25,
	aluifportOut_19,
	dmemaddr26,
	aluifportOut_18,
	dmemaddr27,
	aluifportOut_25,
	dmemaddr28,
	aluifportOut_24,
	dmemaddr29,
	aluifportOut_27,
	dmemaddr30,
	aluifportOut_26,
	dmemaddr31,
	halt_mem,
	dmemstore,
	flush_idex,
	Equal15,
	Equal11,
	Equal0,
	Equal10,
	Equal12,
	Equal20,
	Equal26,
	Equal25,
	Equal13,
	dataScr_ex,
	WideNor0,
	Selector0,
	ALUOP_ex,
	imm_ex,
	ALUScr_ex,
	shamt_ex,
	ALUScr_ex1,
	Regwen_mem,
	regwrite_mem,
	regwrite_mem1,
	regwrite_mem2,
	regwrite_mem3,
	regwrite_mem4,
	rt_ex,
	rt_ex1,
	rt_ex2,
	rt_ex3,
	rt_ex4,
	Regwen_wb,
	regwrite_wb,
	regwrite_wb1,
	regwrite_wb2,
	regwrite_wb3,
	regwrite_wb4,
	dmemload_wb,
	dmemaddr_wb,
	dataScr_wb,
	dataScr_wb1,
	prifpc_mem_1,
	pc_wb,
	Mux622,
	Mux623,
	rdat2_ex,
	prifrs_ex_01,
	prifrs_ex_11,
	prifrs_ex_02,
	prifrs_ex_31,
	prifrs_ex_21,
	prifrs_ex_41,
	opcode_mem,
	opcode_mem1,
	opcode_mem2,
	opcode_mem3,
	opcode_mem4,
	opcode_mem5,
	Mux30,
	Mux301,
	rdat1_ex,
	imm_ex1,
	shamt_ex1,
	dmemload_wb1,
	dmemaddr_wb1,
	prifpc_mem_0,
	pc_wb1,
	Mux632,
	Mux633,
	rdat2_ex1,
	Mux31,
	Mux311,
	rdat1_ex1,
	dmemload_wb2,
	dmemaddr_wb2,
	prifpc_mem_3,
	pc_wb2,
	Mux60,
	Mux601,
	rdat2_ex2,
	imm_ex2,
	shamt_ex2,
	imm_ex3,
	shamt_ex3,
	dmemload_wb3,
	dmemaddr_wb3,
	prifpc_mem_2,
	pc_wb3,
	Mux611,
	Mux612,
	rdat2_ex3,
	dmemload_wb4,
	dmemaddr_wb4,
	prifpc_mem_4,
	pc_wb4,
	Mux59,
	Mux591,
	rdat2_ex4,
	imm_ex4,
	shamt_ex4,
	instr_ex,
	dmemload_wb5,
	imm_wb,
	dmemaddr_wb5,
	pc_wb5,
	Mux321,
	Mux322,
	rdat2_ex5,
	imm_mem,
	imm_wb1,
	dmemload_wb6,
	dmemaddr_wb6,
	pc_wb6,
	Mux331,
	Mux332,
	rdat2_ex6,
	imm_mem1,
	dmemload_wb7,
	imm_wb2,
	dmemaddr_wb7,
	pc_wb7,
	Mux341,
	Mux342,
	rdat2_ex7,
	imm_mem2,
	imm_ex5,
	dmemload_wb8,
	dmemaddr_wb8,
	prifpc_mem_5,
	pc_wb8,
	Mux58,
	Mux581,
	rdat2_ex8,
	imm_ex6,
	dmemload_wb9,
	dmemaddr_wb9,
	prifpc_mem_15,
	pc_wb9,
	Mux48,
	Mux481,
	rdat2_ex9,
	imm_ex7,
	dmemload_wb10,
	dmemaddr_wb10,
	prifpc_mem_14,
	pc_wb10,
	Mux49,
	Mux491,
	rdat2_ex10,
	imm_ex8,
	dmemload_wb11,
	dmemaddr_wb11,
	prifpc_mem_13,
	pc_wb11,
	Mux50,
	Mux501,
	rdat2_ex11,
	imm_ex9,
	dmemload_wb12,
	dmemaddr_wb12,
	prifpc_mem_12,
	pc_wb12,
	Mux51,
	Mux511,
	rdat2_ex12,
	imm_ex10,
	dmemload_wb13,
	dmemaddr_wb13,
	prifpc_mem_11,
	pc_wb13,
	Mux52,
	Mux521,
	rdat2_ex13,
	imm_ex11,
	dmemload_wb14,
	dmemaddr_wb14,
	prifpc_mem_10,
	pc_wb14,
	Mux53,
	Mux531,
	rdat2_ex14,
	imm_ex12,
	dmemload_wb15,
	dmemaddr_wb15,
	prifpc_mem_9,
	pc_wb15,
	Mux54,
	Mux541,
	rdat2_ex15,
	imm_ex13,
	dmemload_wb16,
	dmemaddr_wb16,
	prifpc_mem_6,
	pc_wb16,
	Mux57,
	Mux571,
	rdat2_ex16,
	dmemload_wb17,
	imm_wb3,
	dmemaddr_wb17,
	prifpc_mem_27,
	pc_wb17,
	Mux361,
	Mux362,
	rdat2_ex17,
	imm_mem3,
	dmemload_wb18,
	imm_wb4,
	dmemaddr_wb18,
	prifpc_mem_23,
	pc_wb18,
	Mux401,
	Mux402,
	rdat2_ex18,
	imm_mem4,
	imm_wb5,
	dmemload_wb19,
	dmemaddr_wb19,
	prifpc_mem_18,
	pc_wb19,
	Mux451,
	Mux452,
	rdat2_ex19,
	imm_mem5,
	imm_wb6,
	dmemload_wb20,
	dmemaddr_wb20,
	prifpc_mem_24,
	pc_wb20,
	Mux391,
	Mux392,
	rdat2_ex20,
	imm_mem6,
	imm_wb7,
	dmemload_wb21,
	dmemaddr_wb21,
	prifpc_mem_16,
	pc_wb21,
	Mux471,
	Mux472,
	rdat2_ex21,
	imm_mem7,
	dmemload_wb22,
	imm_wb8,
	dmemaddr_wb22,
	prifpc_mem_19,
	pc_wb22,
	Mux441,
	Mux442,
	rdat2_ex22,
	imm_mem8,
	dmemload_wb23,
	imm_wb9,
	dmemaddr_wb23,
	prifpc_mem_17,
	pc_wb23,
	Mux461,
	Mux462,
	rdat2_ex23,
	imm_mem9,
	dmemload_wb24,
	imm_wb10,
	dmemaddr_wb24,
	prifpc_mem_21,
	pc_wb24,
	Mux421,
	Mux422,
	rdat2_ex24,
	imm_mem10,
	imm_wb11,
	dmemload_wb25,
	dmemaddr_wb25,
	prifpc_mem_20,
	pc_wb25,
	Mux431,
	Mux432,
	rdat2_ex25,
	imm_mem11,
	imm_wb12,
	dmemload_wb26,
	dmemaddr_wb26,
	pc_wb26,
	Mux351,
	Mux352,
	rdat2_ex26,
	imm_mem12,
	imm_wb13,
	dmemload_wb27,
	dmemaddr_wb27,
	prifpc_mem_26,
	pc_wb27,
	Mux371,
	Mux372,
	rdat2_ex27,
	imm_mem13,
	imm_ex14,
	dmemload_wb28,
	dmemaddr_wb28,
	prifpc_mem_8,
	pc_wb28,
	Mux55,
	Mux551,
	rdat2_ex28,
	imm_ex15,
	dmemload_wb29,
	dmemaddr_wb29,
	prifpc_mem_7,
	pc_wb29,
	Mux56,
	Mux561,
	rdat2_ex29,
	imm_wb14,
	dmemload_wb30,
	dmemaddr_wb30,
	prifpc_mem_22,
	pc_wb30,
	Mux411,
	Mux412,
	rdat2_ex30,
	imm_mem14,
	dmemload_wb31,
	imm_wb15,
	dmemaddr_wb31,
	prifpc_mem_25,
	pc_wb31,
	Mux381,
	Mux382,
	rdat2_ex31,
	imm_mem15,
	Equal4,
	ALUOP_ex1,
	Selector2,
	Selector21,
	ALUOP_ex2,
	Mux29,
	Mux291,
	rdat1_ex2,
	Mux27,
	Mux271,
	rdat1_ex3,
	Mux28,
	Mux281,
	rdat1_ex4,
	Mux23,
	Mux231,
	rdat1_ex5,
	Mux24,
	Mux241,
	rdat1_ex6,
	Mux25,
	Mux251,
	rdat1_ex7,
	Mux26,
	Mux261,
	rdat1_ex8,
	Mux15,
	Mux151,
	rdat1_ex9,
	Mux16,
	Mux161,
	rdat1_ex10,
	Mux17,
	Mux171,
	rdat1_ex11,
	Mux18,
	Mux181,
	rdat1_ex12,
	Mux20,
	Mux201,
	rdat1_ex13,
	Mux19,
	Mux191,
	rdat1_ex14,
	Mux21,
	Mux211,
	rdat1_ex15,
	Mux22,
	Mux221,
	rdat1_ex16,
	Mux13,
	Mux131,
	rdat1_ex17,
	Mux14,
	Mux141,
	rdat1_ex18,
	Mux11,
	Mux111,
	rdat1_ex19,
	Mux12,
	Mux121,
	rdat1_ex20,
	Mux9,
	Mux91,
	rdat1_ex21,
	Mux10,
	Mux101,
	rdat1_ex22,
	Mux7,
	Mux71,
	rdat1_ex23,
	Mux8,
	Mux81,
	rdat1_ex24,
	Mux0,
	Mux01,
	rdat1_ex25,
	Mux1,
	Mux110,
	rdat1_ex26,
	Mux2,
	Mux210,
	rdat1_ex27,
	Mux5,
	Mux510,
	rdat1_ex28,
	Mux6,
	Mux64,
	rdat1_ex29,
	Mux3,
	Mux310,
	rdat1_ex30,
	Mux4,
	Mux410,
	rdat1_ex31,
	ALUScr_ex2,
	Selector3,
	ALUOP_ex3,
	aluifportOut_53,
	instr_mem,
	instr_mem1,
	instr_mem2,
	instr_mem3,
	instr_mem4,
	instr_mem5,
	rdat1_mem,
	PCScr_mem,
	pc_bran_mem,
	PCScr_mem1,
	opcode_ex,
	opcode_ex1,
	opcode_ex2,
	opcode_ex3,
	opcode_ex4,
	Equal131,
	memren_ex,
	memwen_ex,
	rdat1_mem1,
	pc_bran_mem1,
	rdat1_mem2,
	pc_bran_mem2,
	rdat1_mem3,
	pc_bran_mem3,
	rdat1_mem4,
	pc_bran_mem4,
	rdat1_mem5,
	pc_bran_mem5,
	rdat1_mem6,
	pc_bran_mem6,
	rdat1_mem7,
	pc_bran_mem7,
	rdat1_mem8,
	pc_bran_mem8,
	instr_mem6,
	rdat1_mem9,
	pc_bran_mem9,
	instr_mem7,
	rdat1_mem10,
	pc_bran_mem10,
	instr_mem8,
	rdat1_mem11,
	pc_bran_mem11,
	instr_mem9,
	rdat1_mem12,
	pc_bran_mem12,
	instr_mem10,
	rdat1_mem13,
	pc_bran_mem13,
	instr_mem11,
	rdat1_mem14,
	pc_bran_mem14,
	instr_mem12,
	rdat1_mem15,
	pc_bran_mem15,
	instr_mem13,
	rdat1_mem16,
	pc_bran_mem16,
	instr_mem14,
	rdat1_mem17,
	pc_bran_mem17,
	instr_mem15,
	rdat1_mem18,
	pc_bran_mem18,
	instr_mem16,
	rdat1_mem19,
	pc_bran_mem19,
	prifpc_mem_151,
	prifpc_mem_291,
	rdat1_mem20,
	pc_bran_mem20,
	prifpc_mem_281,
	rdat1_mem21,
	pc_bran_mem21,
	prifpc_mem_311,
	rdat1_mem22,
	pc_bran_mem22,
	prifpc_mem_301,
	rdat1_mem23,
	pc_bran_mem23,
	instr_mem17,
	rdat1_mem24,
	pc_bran_mem24,
	instr_mem18,
	rdat1_mem25,
	pc_bran_mem25,
	instr_mem19,
	rdat1_mem26,
	pc_bran_mem26,
	instr_mem20,
	rdat1_mem27,
	pc_bran_mem27,
	instr_mem21,
	rdat1_mem28,
	pc_bran_mem28,
	instr_mem22,
	rdat1_mem29,
	pc_bran_mem29,
	instr_mem23,
	rdat1_mem30,
	pc_bran_mem30,
	instr_mem24,
	rdat1_mem31,
	pc_bran_mem31,
	instr_mem25,
	dmemstore1,
	dmemstore2,
	Mux602,
	dmemstore3,
	Mux592,
	dmemstore4,
	Mux582,
	dmemstore5,
	Mux572,
	dmemstore6,
	Mux562,
	dmemstore7,
	Mux552,
	dmemstore8,
	Mux542,
	dmemstore9,
	Mux532,
	dmemstore10,
	Mux522,
	dmemstore11,
	Mux512,
	dmemstore12,
	Mux502,
	dmemstore13,
	Mux492,
	dmemstore14,
	Mux482,
	dmemstore15,
	dmemstore16,
	dmemstore17,
	dmemstore18,
	dmemstore19,
	dmemstore20,
	dmemstore21,
	dmemstore22,
	dmemstore23,
	dmemstore24,
	dmemstore25,
	dmemstore26,
	dmemstore27,
	dmemstore28,
	dmemstore29,
	dmemstore30,
	dmemstore31,
	halt_ex,
	prifhalt_wb,
	ifid_en,
	imemload_id,
	imemload_id1,
	imemload_id2,
	imemload_id3,
	imemload_id4,
	imemload_id5,
	imemload_id6,
	imemload_id7,
	imemload_id8,
	imemload_id9,
	imemload_id10,
	imemload_id11,
	imemload_id12,
	Regwen_ex,
	rd_ex,
	RegDest_ex,
	RegDest_ex1,
	rd_ex1,
	rd_ex2,
	rd_ex3,
	rd_ex4,
	imemload_id13,
	imemload_id14,
	imemload_id15,
	imemload_id16,
	imemload_id17,
	dataScr_mem,
	dataScr_mem1,
	prifpc_mem_110,
	imemload_id18,
	imemload_id19,
	imemload_id20,
	imemload_id21,
	imemload_id22,
	opcode_ex5,
	imemload_id23,
	prifpc_mem_01,
	prifpc_mem_32,
	imemload_id24,
	imemload_id25,
	prifpc_mem_210,
	prifpc_mem_41,
	imemload_id26,
	imemload_id27,
	prifpc_mem_51,
	prifpc_mem_152,
	imemload_id28,
	prifpc_mem_141,
	imemload_id29,
	prifpc_mem_131,
	imemload_id30,
	prifpc_mem_121,
	imemload_id31,
	prifpc_mem_111,
	prifpc_mem_101,
	prifpc_mem_91,
	prifpc_mem_61,
	prifpc_mem_271,
	prifpc_mem_231,
	prifpc_mem_181,
	prifpc_mem_241,
	prifpc_mem_161,
	prifpc_mem_191,
	prifpc_mem_171,
	prifpc_mem_211,
	prifpc_mem_201,
	prifpc_mem_261,
	prifpc_mem_81,
	prifpc_mem_71,
	prifpc_mem_221,
	prifpc_mem_251,
	instr_ex1,
	instr_ex2,
	instr_ex3,
	instr_ex4,
	instr_ex5,
	instr_ex6,
	PCScr_ex,
	pc_ex,
	PCScr_ex1,
	pc_ex1,
	pc_ex2,
	pc_ex3,
	pc_ex4,
	pc_ex5,
	pc_ex6,
	pc_ex7,
	pc_ex8,
	pc_ex9,
	instr_ex7,
	instr_ex8,
	pc_ex10,
	pc_ex11,
	instr_ex9,
	instr_ex10,
	pc_ex12,
	pc_ex13,
	instr_ex11,
	instr_ex12,
	pc_ex14,
	pc_ex15,
	instr_ex13,
	instr_ex14,
	pc_ex16,
	pc_ex17,
	pc_ex18,
	pc_ex19,
	pc_ex20,
	pc_ex21,
	pc_ex22,
	pc_ex23,
	instr_ex15,
	instr_ex16,
	instr_ex17,
	pc_ex24,
	pc_ex25,
	pc_ex26,
	pc_ex27,
	pc_ex28,
	pc_ex29,
	pc_ex30,
	pc_ex31,
	instr_ex18,
	instr_ex19,
	instr_ex20,
	instr_ex21,
	instr_ex22,
	instr_ex23,
	instr_ex24,
	instr_ex25,
	halt_wb,
	dataScr_ex1,
	pc_id,
	pc_id1,
	pc_id2,
	pc_id3,
	pc_id4,
	pc_id5,
	pc_id6,
	pc_id7,
	pc_id8,
	pc_id9,
	pc_id10,
	pc_id11,
	pc_id12,
	pc_id13,
	pc_id14,
	pc_id15,
	pc_id16,
	pc_id17,
	pc_id18,
	pc_id19,
	pc_id20,
	pc_id21,
	pc_id22,
	pc_id23,
	pc_id24,
	pc_id25,
	pc_id26,
	pc_id27,
	pc_id28,
	pc_id29,
	pc_id30,
	pc_id31,
	dataScr_ex2,
	ALUScr_ex3,
	zero_flag_mem,
	devpor,
	devclrn,
	devoe);
input 	prifdmemaddr_1;
input 	pc_1;
input 	prifdmemren;
input 	prifdmemwen;
input 	prifdmemaddr_0;
input 	pc_0;
input 	prifdmemaddr_3;
input 	prifdmemaddr_2;
input 	prifdmemaddr_5;
input 	prifdmemaddr_4;
input 	prifdmemaddr_7;
input 	prifdmemaddr_6;
input 	prifdmemaddr_9;
input 	prifdmemaddr_8;
input 	prifdmemaddr_11;
input 	prifdmemaddr_10;
input 	prifdmemaddr_13;
input 	prifdmemaddr_12;
input 	prifdmemaddr_15;
input 	prifdmemaddr_14;
input 	prifdmemaddr_23;
input 	prifdmemaddr_22;
input 	prifdmemaddr_21;
input 	prifdmemaddr_29;
input 	prifdmemaddr_28;
input 	prifdmemaddr_31;
input 	prifdmemaddr_30;
input 	prifdmemaddr_20;
input 	prifdmemaddr_17;
input 	prifdmemaddr_16;
input 	prifdmemaddr_19;
input 	prifdmemaddr_18;
input 	prifdmemaddr_25;
input 	prifdmemaddr_24;
input 	prifdmemaddr_27;
input 	prifdmemaddr_26;
input 	prifhalt_mem;
input 	prifdmemstore_0;
input 	prifimm_ex_1;
input 	prifALUScr_ex_1;
input 	prifshamt_ex_1;
input 	prifALUScr_ex_0;
input 	prifRegwen_mem;
input 	prifregwrite_mem_4;
input 	prifregwrite_mem_0;
input 	prifregwrite_mem_1;
input 	prifregwrite_mem_2;
input 	prifregwrite_mem_3;
input 	prifrt_ex_1;
input 	prifrt_ex_0;
input 	prifrt_ex_3;
input 	prifrt_ex_2;
input 	prifrt_ex_4;
input 	prifrdat2_ex_1;
input 	prifopcode_mem_1;
input 	prifopcode_mem_0;
input 	prifopcode_mem_2;
input 	prifopcode_mem_3;
input 	prifopcode_mem_5;
input 	prifopcode_mem_4;
input 	prifrdat1_ex_1;
input 	prifimm_ex_0;
input 	prifshamt_ex_0;
input 	prifrdat2_ex_0;
input 	prifrdat1_ex_0;
input 	prifrdat2_ex_3;
input 	prifimm_ex_3;
input 	prifshamt_ex_3;
input 	prifimm_ex_2;
input 	prifshamt_ex_2;
input 	prifrdat2_ex_2;
input 	prifrdat2_ex_4;
input 	prifimm_ex_4;
input 	prifshamt_ex_4;
input 	prifinstr_ex_15;
input 	prifrdat2_ex_31;
input 	prifimm_mem_15;
input 	prifrdat2_ex_30;
input 	prifimm_mem_14;
input 	prifrdat2_ex_29;
input 	prifimm_mem_13;
input 	prifimm_ex_5;
input 	prifrdat2_ex_5;
input 	prifimm_ex_15;
input 	prifrdat2_ex_15;
input 	prifimm_ex_14;
input 	prifrdat2_ex_14;
input 	prifimm_ex_13;
input 	prifrdat2_ex_13;
input 	prifimm_ex_12;
input 	prifrdat2_ex_12;
input 	prifimm_ex_11;
input 	prifrdat2_ex_11;
input 	prifimm_ex_10;
input 	prifrdat2_ex_10;
input 	prifimm_ex_9;
input 	prifrdat2_ex_9;
input 	prifimm_ex_6;
input 	prifrdat2_ex_6;
input 	prifrdat2_ex_27;
input 	prifimm_mem_11;
input 	prifrdat2_ex_23;
input 	prifimm_mem_7;
input 	prifrdat2_ex_18;
input 	prifimm_mem_2;
input 	prifrdat2_ex_24;
input 	prifimm_mem_8;
input 	prifrdat2_ex_16;
input 	prifimm_mem_0;
input 	prifrdat2_ex_19;
input 	prifimm_mem_3;
input 	prifrdat2_ex_17;
input 	prifimm_mem_1;
input 	prifrdat2_ex_21;
input 	prifimm_mem_5;
input 	prifrdat2_ex_20;
input 	prifimm_mem_4;
input 	prifrdat2_ex_28;
input 	prifimm_mem_12;
input 	prifrdat2_ex_26;
input 	prifimm_mem_10;
input 	prifimm_ex_8;
input 	prifrdat2_ex_8;
input 	prifimm_ex_7;
input 	prifrdat2_ex_7;
input 	prifrdat2_ex_22;
input 	prifimm_mem_6;
input 	prifrdat2_ex_25;
input 	prifimm_mem_9;
input 	prifrdat1_ex_2;
input 	prifrdat1_ex_4;
input 	prifrdat1_ex_3;
input 	prifrdat1_ex_8;
input 	prifrdat1_ex_7;
input 	prifrdat1_ex_6;
input 	prifrdat1_ex_5;
input 	prifrdat1_ex_16;
input 	prifrdat1_ex_15;
input 	prifrdat1_ex_14;
input 	prifrdat1_ex_13;
input 	prifrdat1_ex_11;
input 	prifrdat1_ex_12;
input 	prifrdat1_ex_10;
input 	prifrdat1_ex_9;
input 	prifrdat1_ex_18;
input 	prifrdat1_ex_17;
input 	prifrdat1_ex_20;
input 	prifrdat1_ex_19;
input 	prifrdat1_ex_22;
input 	prifrdat1_ex_21;
input 	prifrdat1_ex_24;
input 	prifrdat1_ex_23;
input 	prifrdat1_ex_31;
input 	prifrdat1_ex_30;
input 	prifrdat1_ex_29;
input 	prifrdat1_ex_26;
input 	prifrdat1_ex_25;
input 	prifrdat1_ex_28;
input 	prifrdat1_ex_27;
input 	prifzero_flag_mem;
input 	prifinstr_mem_3;
input 	prifinstr_mem_5;
input 	prifinstr_mem_4;
input 	prifinstr_mem_2;
input 	prifinstr_mem_1;
input 	prifinstr_mem_0;
input 	prifrdat1_mem_1;
input 	prifPCScr_mem_0;
input 	prifpc_bran_mem_1;
input 	prifPCScr_mem_1;
input 	prifopcode_ex_5;
input 	prifopcode_ex_0;
input 	prifopcode_ex_1;
input 	prifopcode_ex_2;
input 	prifopcode_ex_4;
input 	prifmemren_ex;
input 	prifmemwen_ex;
input 	prifrdat1_mem_0;
input 	prifpc_bran_mem_0;
input 	prifrdat1_mem_3;
input 	prifpc_bran_mem_3;
input 	prifrdat1_mem_2;
input 	prifpc_bran_mem_2;
input 	prifrdat1_mem_5;
input 	prifpc_bran_mem_5;
input 	prifrdat1_mem_4;
input 	prifpc_bran_mem_4;
input 	prifrdat1_mem_7;
input 	prifpc_bran_mem_7;
input 	prifrdat1_mem_6;
input 	prifpc_bran_mem_6;
input 	prifrdat1_mem_9;
input 	prifpc_bran_mem_9;
input 	prifinstr_mem_7;
input 	prifrdat1_mem_8;
input 	prifpc_bran_mem_8;
input 	prifinstr_mem_6;
input 	prifrdat1_mem_11;
input 	prifpc_bran_mem_11;
input 	prifinstr_mem_9;
input 	prifrdat1_mem_10;
input 	prifpc_bran_mem_10;
input 	prifinstr_mem_8;
input 	prifrdat1_mem_13;
input 	prifpc_bran_mem_13;
input 	prifinstr_mem_11;
input 	prifrdat1_mem_12;
input 	prifpc_bran_mem_12;
input 	prifinstr_mem_10;
input 	prifrdat1_mem_15;
input 	prifpc_bran_mem_15;
input 	prifinstr_mem_13;
input 	prifrdat1_mem_14;
input 	prifpc_bran_mem_14;
input 	prifinstr_mem_12;
input 	prifrdat1_mem_23;
input 	prifpc_bran_mem_23;
input 	prifinstr_mem_21;
input 	prifrdat1_mem_22;
input 	prifpc_bran_mem_22;
input 	prifinstr_mem_20;
input 	prifrdat1_mem_21;
input 	prifpc_bran_mem_21;
input 	prifinstr_mem_19;
input 	prifrdat1_mem_29;
input 	prifpc_bran_mem_29;
input 	prifrdat1_mem_28;
input 	prifpc_bran_mem_28;
input 	prifrdat1_mem_31;
input 	prifpc_bran_mem_31;
input 	prifrdat1_mem_30;
input 	prifpc_bran_mem_30;
input 	prifrdat1_mem_20;
input 	prifpc_bran_mem_20;
input 	prifinstr_mem_18;
input 	prifrdat1_mem_17;
input 	prifpc_bran_mem_17;
input 	prifinstr_mem_15;
input 	prifrdat1_mem_16;
input 	prifpc_bran_mem_16;
input 	prifinstr_mem_14;
input 	prifrdat1_mem_19;
input 	prifpc_bran_mem_19;
input 	prifinstr_mem_17;
input 	prifrdat1_mem_18;
input 	prifpc_bran_mem_18;
input 	prifinstr_mem_16;
input 	prifrdat1_mem_25;
input 	prifpc_bran_mem_25;
input 	prifinstr_mem_23;
input 	prifrdat1_mem_24;
input 	prifpc_bran_mem_24;
input 	prifinstr_mem_22;
input 	prifrdat1_mem_27;
input 	prifpc_bran_mem_27;
input 	prifinstr_mem_25;
input 	prifrdat1_mem_26;
input 	prifpc_bran_mem_26;
input 	prifinstr_mem_24;
input 	prifdmemstore_1;
input 	prifdmemstore_2;
input 	prifdmemstore_3;
input 	prifdmemstore_4;
input 	prifdmemstore_5;
input 	prifdmemstore_6;
input 	prifdmemstore_7;
input 	prifdmemstore_8;
input 	prifdmemstore_9;
input 	prifdmemstore_10;
input 	prifdmemstore_11;
input 	prifdmemstore_12;
input 	prifdmemstore_13;
input 	prifdmemstore_14;
input 	prifdmemstore_15;
input 	prifdmemstore_16;
input 	prifdmemstore_17;
input 	prifdmemstore_18;
input 	prifdmemstore_19;
input 	prifdmemstore_20;
input 	prifdmemstore_21;
input 	prifdmemstore_22;
input 	prifdmemstore_23;
input 	prifdmemstore_24;
input 	prifdmemstore_25;
input 	prifdmemstore_26;
input 	prifdmemstore_27;
input 	prifdmemstore_28;
input 	prifdmemstore_29;
input 	prifdmemstore_30;
input 	prifdmemstore_31;
input 	prifhalt_ex;
input 	prifimemload_id_31;
input 	prifimemload_id_30;
input 	prifimemload_id_29;
input 	prifimemload_id_27;
input 	prifimemload_id_26;
input 	prifimemload_id_28;
input 	prifimemload_id_3;
input 	prifimemload_id_1;
input 	prifimemload_id_5;
input 	prifimemload_id_4;
input 	prifimemload_id_2;
input 	prifimemload_id_0;
input 	prifimemload_id_7;
input 	prifRegwen_ex;
input 	prifrd_ex_4;
input 	prifRegDest_ex_1;
input 	prifRegDest_ex_0;
input 	prifrd_ex_0;
input 	prifrd_ex_1;
input 	prifrd_ex_2;
input 	prifrd_ex_3;
input 	prifimemload_id_17;
input 	prifimemload_id_16;
input 	prifimemload_id_19;
input 	prifimemload_id_18;
input 	prifimemload_id_20;
input 	prifdataScr_mem_0;
input 	prifdataScr_mem_1;
input 	prifimemload_id_22;
input 	prifimemload_id_21;
input 	prifimemload_id_24;
input 	prifimemload_id_23;
input 	prifimemload_id_25;
input 	prifopcode_ex_3;
input 	prifimemload_id_6;
input 	prifimemload_id_9;
input 	prifimemload_id_8;
input 	prifimemload_id_10;
input 	prifimemload_id_15;
input 	prifimemload_id_14;
input 	prifimemload_id_13;
input 	prifimemload_id_12;
input 	prifimemload_id_11;
input 	prifinstr_ex_3;
input 	prifinstr_ex_5;
input 	prifinstr_ex_4;
input 	prifinstr_ex_2;
input 	prifinstr_ex_1;
input 	prifinstr_ex_0;
input 	prifPCScr_ex_0;
input 	prifpc_ex_1;
input 	prifPCScr_ex_1;
input 	prifpc_ex_0;
input 	prifpc_ex_3;
input 	prifpc_ex_2;
input 	Add0;
input 	Add01;
input 	prifpc_ex_5;
input 	prifpc_ex_4;
input 	Add02;
input 	Add03;
input 	prifpc_ex_7;
input 	prifpc_ex_6;
input 	Add04;
input 	Add05;
input 	prifpc_ex_9;
input 	prifpc_ex_8;
input 	Add06;
input 	Add07;
input 	prifinstr_ex_7;
input 	prifinstr_ex_6;
input 	prifpc_ex_11;
input 	prifpc_ex_10;
input 	Add08;
input 	Add09;
input 	prifinstr_ex_9;
input 	prifinstr_ex_8;
input 	prifpc_ex_13;
input 	prifpc_ex_12;
input 	Add010;
input 	Add011;
input 	prifinstr_ex_11;
input 	prifinstr_ex_10;
input 	prifpc_ex_15;
input 	prifpc_ex_14;
input 	Add012;
input 	Add013;
input 	prifinstr_ex_13;
input 	prifinstr_ex_12;
input 	prifpc_ex_23;
input 	prifpc_ex_22;
input 	prifpc_ex_21;
input 	prifpc_ex_20;
input 	prifpc_ex_19;
input 	prifpc_ex_18;
input 	prifpc_ex_17;
input 	prifpc_ex_16;
input 	Add014;
input 	Add015;
input 	Add016;
input 	Add017;
input 	Add018;
input 	Add019;
input 	Add020;
input 	Add021;
input 	prifinstr_ex_21;
input 	prifinstr_ex_20;
input 	prifinstr_ex_19;
input 	prifpc_ex_29;
input 	prifpc_ex_28;
input 	prifpc_ex_27;
input 	prifpc_ex_26;
input 	prifpc_ex_25;
input 	prifpc_ex_24;
input 	Add022;
input 	Add023;
input 	Add024;
input 	Add025;
input 	Add026;
input 	Add027;
input 	prifpc_ex_31;
input 	prifpc_ex_30;
input 	Add028;
input 	Add029;
input 	prifinstr_ex_18;
input 	prifinstr_ex_14;
input 	prifinstr_ex_17;
input 	prifinstr_ex_16;
input 	prifinstr_ex_23;
input 	prifinstr_ex_22;
input 	prifinstr_ex_25;
input 	prifinstr_ex_24;
input 	prifdataScr_ex_0;
input 	prifdataScr_ex_1;
input 	prifpc_id_1;
input 	prifpc_id_0;
input 	prifpc_id_3;
input 	prifpc_id_2;
input 	prifpc_id_5;
input 	prifpc_id_4;
input 	prifpc_id_7;
input 	prifpc_id_6;
input 	prifpc_id_9;
input 	prifpc_id_8;
input 	prifpc_id_11;
input 	prifpc_id_10;
input 	prifpc_id_13;
input 	prifpc_id_12;
input 	prifpc_id_15;
input 	prifpc_id_14;
input 	prifpc_id_23;
input 	prifpc_id_22;
input 	prifpc_id_21;
input 	prifpc_id_20;
input 	prifpc_id_19;
input 	prifpc_id_18;
input 	prifpc_id_17;
input 	prifpc_id_16;
input 	prifpc_id_29;
input 	prifpc_id_28;
input 	prifpc_id_27;
input 	prifpc_id_26;
input 	prifpc_id_25;
input 	prifpc_id_24;
input 	prifpc_id_31;
input 	prifpc_id_30;
input 	Add2;
input 	Add21;
input 	Add22;
input 	Add23;
input 	Add24;
input 	Add25;
input 	Add26;
input 	Add27;
input 	Add28;
input 	Add29;
input 	Add210;
input 	Add211;
input 	Add212;
input 	Add213;
input 	Add214;
input 	Add215;
input 	Add216;
input 	Add217;
input 	Add218;
input 	Add219;
input 	Add220;
input 	Add221;
input 	Add222;
input 	Add223;
input 	Add224;
input 	Add225;
input 	Add226;
input 	Add227;
input 	Add228;
input 	pc_2;
input 	always1;
input 	ramiframload_0;
input 	ramiframload_1;
input 	ramiframload_2;
input 	ramiframload_3;
input 	ramiframload_4;
input 	ramiframload_5;
input 	ramiframload_6;
input 	ramiframload_7;
input 	ramiframload_8;
input 	ramiframload_9;
input 	ramiframload_10;
input 	ramiframload_11;
input 	ramiframload_12;
input 	ramiframload_13;
input 	ramiframload_14;
input 	ramiframload_15;
input 	ramiframload_16;
input 	ramiframload_17;
input 	ramiframload_18;
input 	ramiframload_19;
input 	ramiframload_20;
input 	ramiframload_21;
input 	ramiframload_22;
input 	ramiframload_23;
input 	ramiframload_24;
input 	ramiframload_25;
input 	ramiframload_26;
input 	ramiframload_27;
input 	ramiframload_28;
input 	ramiframload_29;
input 	ramiframload_30;
input 	ramiframload_31;
input 	prifALUOP_ex_3;
input 	prifRegwen_wb;
input 	prifregwrite_wb_2;
input 	prifregwrite_wb_0;
input 	prifregwrite_wb_1;
input 	prifregwrite_wb_4;
input 	prifregwrite_wb_3;
input 	Mux62;
input 	prifdmemload_wb_1;
input 	prifdmemaddr_wb_1;
input 	prifdataScr_wb_0;
input 	prifdataScr_wb_1;
input 	prifpc_wb_1;
input 	Mux621;
input 	prifrs_ex_1;
input 	prifrs_ex_0;
input 	prifrs_ex_3;
input 	prifrs_ex_2;
input 	prifrs_ex_4;
input 	Mux63;
input 	prifdmemload_wb_0;
input 	prifdmemaddr_wb_0;
input 	prifpc_wb_0;
input 	Mux631;
input 	prifdmemload_wb_3;
input 	prifdmemaddr_wb_3;
input 	prifpc_wb_3;
input 	prifdmemload_wb_2;
input 	prifdmemaddr_wb_2;
input 	prifpc_wb_2;
input 	Mux61;
input 	prifdmemload_wb_4;
input 	prifdmemaddr_wb_4;
input 	prifpc_wb_4;
input 	prifdmemload_wb_31;
input 	prifimm_wb_15;
input 	prifdmemaddr_wb_31;
input 	prifpc_wb_31;
input 	Mux32;
input 	prifimm_wb_14;
input 	prifdmemload_wb_30;
input 	prifdmemaddr_wb_30;
input 	prifpc_wb_30;
input 	Mux33;
input 	prifdmemload_wb_29;
input 	prifimm_wb_13;
input 	prifdmemaddr_wb_29;
input 	prifpc_wb_29;
input 	Mux34;
input 	prifdmemload_wb_5;
input 	prifdmemaddr_wb_5;
input 	prifpc_wb_5;
input 	prifdmemload_wb_15;
input 	prifdmemaddr_wb_15;
input 	prifpc_wb_15;
input 	prifdmemload_wb_14;
input 	prifdmemaddr_wb_14;
input 	prifpc_wb_14;
input 	prifdmemload_wb_13;
input 	prifdmemaddr_wb_13;
input 	prifpc_wb_13;
input 	prifdmemload_wb_12;
input 	prifdmemaddr_wb_12;
input 	prifpc_wb_12;
input 	prifdmemload_wb_11;
input 	prifdmemaddr_wb_11;
input 	prifpc_wb_11;
input 	prifdmemload_wb_10;
input 	prifdmemaddr_wb_10;
input 	prifpc_wb_10;
input 	prifdmemload_wb_9;
input 	prifdmemaddr_wb_9;
input 	prifpc_wb_9;
input 	prifdmemload_wb_6;
input 	prifdmemaddr_wb_6;
input 	prifpc_wb_6;
input 	prifdmemload_wb_27;
input 	prifimm_wb_11;
input 	prifdmemaddr_wb_27;
input 	prifpc_wb_27;
input 	Mux36;
input 	prifdmemload_wb_23;
input 	prifimm_wb_7;
input 	prifdmemaddr_wb_23;
input 	prifpc_wb_23;
input 	Mux40;
input 	prifimm_wb_2;
input 	prifdmemload_wb_18;
input 	prifdmemaddr_wb_18;
input 	prifpc_wb_18;
input 	Mux45;
input 	prifimm_wb_8;
input 	prifdmemload_wb_24;
input 	prifdmemaddr_wb_24;
input 	prifpc_wb_24;
input 	Mux39;
input 	prifimm_wb_0;
input 	prifdmemload_wb_16;
input 	prifdmemaddr_wb_16;
input 	prifpc_wb_16;
input 	Mux47;
input 	prifdmemload_wb_19;
input 	prifimm_wb_3;
input 	prifdmemaddr_wb_19;
input 	prifpc_wb_19;
input 	Mux44;
input 	prifdmemload_wb_17;
input 	prifimm_wb_1;
input 	prifdmemaddr_wb_17;
input 	prifpc_wb_17;
input 	Mux46;
input 	prifdmemload_wb_21;
input 	prifimm_wb_5;
input 	prifdmemaddr_wb_21;
input 	prifpc_wb_21;
input 	Mux42;
input 	prifimm_wb_4;
input 	prifdmemload_wb_20;
input 	prifdmemaddr_wb_20;
input 	prifpc_wb_20;
input 	Mux43;
input 	prifimm_wb_12;
input 	prifdmemload_wb_28;
input 	prifdmemaddr_wb_28;
input 	prifpc_wb_28;
input 	Mux35;
input 	prifimm_wb_10;
input 	prifdmemload_wb_26;
input 	prifdmemaddr_wb_26;
input 	prifpc_wb_26;
input 	Mux37;
input 	prifdmemload_wb_8;
input 	prifdmemaddr_wb_8;
input 	prifpc_wb_8;
input 	prifdmemload_wb_7;
input 	prifdmemaddr_wb_7;
input 	prifpc_wb_7;
input 	prifimm_wb_6;
input 	prifdmemload_wb_22;
input 	prifdmemaddr_wb_22;
input 	prifpc_wb_22;
input 	Mux41;
input 	prifdmemload_wb_25;
input 	prifimm_wb_9;
input 	prifdmemaddr_wb_25;
input 	prifpc_wb_25;
input 	Mux38;
input 	prifALUOP_ex_2;
input 	prifALUOP_ex_1;
input 	prifALUOP_ex_0;
input 	aluifportOut_1;
input 	exmem_en;
output 	dmemaddr;
input 	ccifiwait_0;
output 	dmemren;
output 	dmemwen;
input 	aluifportOut_0;
output 	dmemaddr1;
input 	aluifportOut_3;
input 	aluifportOut_5;
input 	aluifportOut_2;
input 	aluifportOut_31;
input 	aluifportOut_32;
output 	dmemaddr2;
input 	aluifportOut_21;
output 	dmemaddr3;
input 	aluifportOut_51;
input 	aluifportOut_52;
output 	dmemaddr4;
input 	aluifportOut_4;
output 	dmemaddr5;
input 	aluifportOut_7;
output 	dmemaddr6;
input 	aluifportOut_6;
output 	dmemaddr7;
input 	aluifportOut_9;
output 	dmemaddr8;
input 	aluifportOut_8;
output 	dmemaddr9;
input 	aluifportOut_11;
output 	dmemaddr10;
input 	aluifportOut_10;
output 	dmemaddr11;
input 	aluifportOut_13;
output 	dmemaddr12;
input 	aluifportOut_12;
output 	dmemaddr13;
input 	aluifportOut_15;
output 	dmemaddr14;
input 	aluifportOut_14;
output 	dmemaddr15;
input 	aluifportOut_23;
output 	dmemaddr16;
input 	aluifportOut_22;
output 	dmemaddr17;
input 	aluifportOut_211;
output 	dmemaddr18;
input 	aluifportOut_29;
output 	dmemaddr19;
input 	prifpc_mem_29;
input 	aluifportOut_28;
output 	dmemaddr20;
input 	prifpc_mem_28;
input 	aluifneg_flag;
output 	dmemaddr21;
input 	prifpc_mem_31;
input 	aluifportOut_30;
output 	dmemaddr22;
input 	prifpc_mem_30;
input 	aluifportOut_20;
output 	dmemaddr23;
input 	aluifportOut_17;
output 	dmemaddr24;
input 	aluifportOut_16;
output 	dmemaddr25;
input 	aluifportOut_19;
output 	dmemaddr26;
input 	aluifportOut_18;
output 	dmemaddr27;
input 	aluifportOut_25;
output 	dmemaddr28;
input 	aluifportOut_24;
output 	dmemaddr29;
input 	aluifportOut_27;
output 	dmemaddr30;
input 	aluifportOut_26;
output 	dmemaddr31;
output 	halt_mem;
output 	dmemstore;
input 	flush_idex;
input 	Equal15;
input 	Equal11;
input 	Equal0;
input 	Equal10;
input 	Equal12;
input 	Equal20;
input 	Equal26;
input 	Equal25;
input 	Equal13;
output 	dataScr_ex;
input 	WideNor0;
input 	Selector0;
output 	ALUOP_ex;
output 	imm_ex;
output 	ALUScr_ex;
output 	shamt_ex;
output 	ALUScr_ex1;
output 	Regwen_mem;
output 	regwrite_mem;
output 	regwrite_mem1;
output 	regwrite_mem2;
output 	regwrite_mem3;
output 	regwrite_mem4;
output 	rt_ex;
output 	rt_ex1;
output 	rt_ex2;
output 	rt_ex3;
output 	rt_ex4;
output 	Regwen_wb;
output 	regwrite_wb;
output 	regwrite_wb1;
output 	regwrite_wb2;
output 	regwrite_wb3;
output 	regwrite_wb4;
output 	dmemload_wb;
output 	dmemaddr_wb;
output 	dataScr_wb;
output 	dataScr_wb1;
input 	prifpc_mem_1;
output 	pc_wb;
input 	Mux622;
input 	Mux623;
output 	rdat2_ex;
input 	prifrs_ex_01;
output 	prifrs_ex_11;
output 	prifrs_ex_02;
output 	prifrs_ex_31;
output 	prifrs_ex_21;
output 	prifrs_ex_41;
output 	opcode_mem;
output 	opcode_mem1;
output 	opcode_mem2;
output 	opcode_mem3;
output 	opcode_mem4;
output 	opcode_mem5;
input 	Mux30;
input 	Mux301;
output 	rdat1_ex;
output 	imm_ex1;
output 	shamt_ex1;
output 	dmemload_wb1;
output 	dmemaddr_wb1;
input 	prifpc_mem_0;
output 	pc_wb1;
input 	Mux632;
input 	Mux633;
output 	rdat2_ex1;
input 	Mux31;
input 	Mux311;
output 	rdat1_ex1;
output 	dmemload_wb2;
output 	dmemaddr_wb2;
input 	prifpc_mem_3;
output 	pc_wb2;
input 	Mux60;
input 	Mux601;
output 	rdat2_ex2;
output 	imm_ex2;
output 	shamt_ex2;
output 	imm_ex3;
output 	shamt_ex3;
output 	dmemload_wb3;
output 	dmemaddr_wb3;
input 	prifpc_mem_2;
output 	pc_wb3;
input 	Mux611;
input 	Mux612;
output 	rdat2_ex3;
output 	dmemload_wb4;
output 	dmemaddr_wb4;
input 	prifpc_mem_4;
output 	pc_wb4;
input 	Mux59;
input 	Mux591;
output 	rdat2_ex4;
output 	imm_ex4;
output 	shamt_ex4;
output 	instr_ex;
output 	dmemload_wb5;
output 	imm_wb;
output 	dmemaddr_wb5;
output 	pc_wb5;
input 	Mux321;
input 	Mux322;
output 	rdat2_ex5;
output 	imm_mem;
output 	imm_wb1;
output 	dmemload_wb6;
output 	dmemaddr_wb6;
output 	pc_wb6;
input 	Mux331;
input 	Mux332;
output 	rdat2_ex6;
output 	imm_mem1;
output 	dmemload_wb7;
output 	imm_wb2;
output 	dmemaddr_wb7;
output 	pc_wb7;
input 	Mux341;
input 	Mux342;
output 	rdat2_ex7;
output 	imm_mem2;
output 	imm_ex5;
output 	dmemload_wb8;
output 	dmemaddr_wb8;
input 	prifpc_mem_5;
output 	pc_wb8;
input 	Mux58;
input 	Mux581;
output 	rdat2_ex8;
output 	imm_ex6;
output 	dmemload_wb9;
output 	dmemaddr_wb9;
input 	prifpc_mem_15;
output 	pc_wb9;
input 	Mux48;
input 	Mux481;
output 	rdat2_ex9;
output 	imm_ex7;
output 	dmemload_wb10;
output 	dmemaddr_wb10;
input 	prifpc_mem_14;
output 	pc_wb10;
input 	Mux49;
input 	Mux491;
output 	rdat2_ex10;
output 	imm_ex8;
output 	dmemload_wb11;
output 	dmemaddr_wb11;
input 	prifpc_mem_13;
output 	pc_wb11;
input 	Mux50;
input 	Mux501;
output 	rdat2_ex11;
output 	imm_ex9;
output 	dmemload_wb12;
output 	dmemaddr_wb12;
input 	prifpc_mem_12;
output 	pc_wb12;
input 	Mux51;
input 	Mux511;
output 	rdat2_ex12;
output 	imm_ex10;
output 	dmemload_wb13;
output 	dmemaddr_wb13;
input 	prifpc_mem_11;
output 	pc_wb13;
input 	Mux52;
input 	Mux521;
output 	rdat2_ex13;
output 	imm_ex11;
output 	dmemload_wb14;
output 	dmemaddr_wb14;
input 	prifpc_mem_10;
output 	pc_wb14;
input 	Mux53;
input 	Mux531;
output 	rdat2_ex14;
output 	imm_ex12;
output 	dmemload_wb15;
output 	dmemaddr_wb15;
input 	prifpc_mem_9;
output 	pc_wb15;
input 	Mux54;
input 	Mux541;
output 	rdat2_ex15;
output 	imm_ex13;
output 	dmemload_wb16;
output 	dmemaddr_wb16;
input 	prifpc_mem_6;
output 	pc_wb16;
input 	Mux57;
input 	Mux571;
output 	rdat2_ex16;
output 	dmemload_wb17;
output 	imm_wb3;
output 	dmemaddr_wb17;
input 	prifpc_mem_27;
output 	pc_wb17;
input 	Mux361;
input 	Mux362;
output 	rdat2_ex17;
output 	imm_mem3;
output 	dmemload_wb18;
output 	imm_wb4;
output 	dmemaddr_wb18;
input 	prifpc_mem_23;
output 	pc_wb18;
input 	Mux401;
input 	Mux402;
output 	rdat2_ex18;
output 	imm_mem4;
output 	imm_wb5;
output 	dmemload_wb19;
output 	dmemaddr_wb19;
input 	prifpc_mem_18;
output 	pc_wb19;
input 	Mux451;
input 	Mux452;
output 	rdat2_ex19;
output 	imm_mem5;
output 	imm_wb6;
output 	dmemload_wb20;
output 	dmemaddr_wb20;
input 	prifpc_mem_24;
output 	pc_wb20;
input 	Mux391;
input 	Mux392;
output 	rdat2_ex20;
output 	imm_mem6;
output 	imm_wb7;
output 	dmemload_wb21;
output 	dmemaddr_wb21;
input 	prifpc_mem_16;
output 	pc_wb21;
input 	Mux471;
input 	Mux472;
output 	rdat2_ex21;
output 	imm_mem7;
output 	dmemload_wb22;
output 	imm_wb8;
output 	dmemaddr_wb22;
input 	prifpc_mem_19;
output 	pc_wb22;
input 	Mux441;
input 	Mux442;
output 	rdat2_ex22;
output 	imm_mem8;
output 	dmemload_wb23;
output 	imm_wb9;
output 	dmemaddr_wb23;
input 	prifpc_mem_17;
output 	pc_wb23;
input 	Mux461;
input 	Mux462;
output 	rdat2_ex23;
output 	imm_mem9;
output 	dmemload_wb24;
output 	imm_wb10;
output 	dmemaddr_wb24;
input 	prifpc_mem_21;
output 	pc_wb24;
input 	Mux421;
input 	Mux422;
output 	rdat2_ex24;
output 	imm_mem10;
output 	imm_wb11;
output 	dmemload_wb25;
output 	dmemaddr_wb25;
input 	prifpc_mem_20;
output 	pc_wb25;
input 	Mux431;
input 	Mux432;
output 	rdat2_ex25;
output 	imm_mem11;
output 	imm_wb12;
output 	dmemload_wb26;
output 	dmemaddr_wb26;
output 	pc_wb26;
input 	Mux351;
input 	Mux352;
output 	rdat2_ex26;
output 	imm_mem12;
output 	imm_wb13;
output 	dmemload_wb27;
output 	dmemaddr_wb27;
input 	prifpc_mem_26;
output 	pc_wb27;
input 	Mux371;
input 	Mux372;
output 	rdat2_ex27;
output 	imm_mem13;
output 	imm_ex14;
output 	dmemload_wb28;
output 	dmemaddr_wb28;
input 	prifpc_mem_8;
output 	pc_wb28;
input 	Mux55;
input 	Mux551;
output 	rdat2_ex28;
output 	imm_ex15;
output 	dmemload_wb29;
output 	dmemaddr_wb29;
input 	prifpc_mem_7;
output 	pc_wb29;
input 	Mux56;
input 	Mux561;
output 	rdat2_ex29;
output 	imm_wb14;
output 	dmemload_wb30;
output 	dmemaddr_wb30;
input 	prifpc_mem_22;
output 	pc_wb30;
input 	Mux411;
input 	Mux412;
output 	rdat2_ex30;
output 	imm_mem14;
output 	dmemload_wb31;
output 	imm_wb15;
output 	dmemaddr_wb31;
input 	prifpc_mem_25;
output 	pc_wb31;
input 	Mux381;
input 	Mux382;
output 	rdat2_ex31;
output 	imm_mem15;
input 	Equal4;
output 	ALUOP_ex1;
input 	Selector2;
input 	Selector21;
output 	ALUOP_ex2;
input 	Mux29;
input 	Mux291;
output 	rdat1_ex2;
input 	Mux27;
input 	Mux271;
output 	rdat1_ex3;
input 	Mux28;
input 	Mux281;
output 	rdat1_ex4;
input 	Mux23;
input 	Mux231;
output 	rdat1_ex5;
input 	Mux24;
input 	Mux241;
output 	rdat1_ex6;
input 	Mux25;
input 	Mux251;
output 	rdat1_ex7;
input 	Mux26;
input 	Mux261;
output 	rdat1_ex8;
input 	Mux15;
input 	Mux151;
output 	rdat1_ex9;
input 	Mux16;
input 	Mux161;
output 	rdat1_ex10;
input 	Mux17;
input 	Mux171;
output 	rdat1_ex11;
input 	Mux18;
input 	Mux181;
output 	rdat1_ex12;
input 	Mux20;
input 	Mux201;
output 	rdat1_ex13;
input 	Mux19;
input 	Mux191;
output 	rdat1_ex14;
input 	Mux21;
input 	Mux211;
output 	rdat1_ex15;
input 	Mux22;
input 	Mux221;
output 	rdat1_ex16;
input 	Mux13;
input 	Mux131;
output 	rdat1_ex17;
input 	Mux14;
input 	Mux141;
output 	rdat1_ex18;
input 	Mux11;
input 	Mux111;
output 	rdat1_ex19;
input 	Mux12;
input 	Mux121;
output 	rdat1_ex20;
input 	Mux9;
input 	Mux91;
output 	rdat1_ex21;
input 	Mux10;
input 	Mux101;
output 	rdat1_ex22;
input 	Mux7;
input 	Mux71;
output 	rdat1_ex23;
input 	Mux8;
input 	Mux81;
output 	rdat1_ex24;
input 	Mux0;
input 	Mux01;
output 	rdat1_ex25;
input 	Mux1;
input 	Mux110;
output 	rdat1_ex26;
input 	Mux2;
input 	Mux210;
output 	rdat1_ex27;
input 	Mux5;
input 	Mux510;
output 	rdat1_ex28;
input 	Mux6;
input 	Mux64;
output 	rdat1_ex29;
input 	Mux3;
input 	Mux310;
output 	rdat1_ex30;
input 	Mux4;
input 	Mux410;
output 	rdat1_ex31;
output 	ALUScr_ex2;
input 	Selector3;
output 	ALUOP_ex3;
input 	aluifportOut_53;
output 	instr_mem;
output 	instr_mem1;
output 	instr_mem2;
output 	instr_mem3;
output 	instr_mem4;
output 	instr_mem5;
output 	rdat1_mem;
output 	PCScr_mem;
output 	pc_bran_mem;
output 	PCScr_mem1;
output 	opcode_ex;
output 	opcode_ex1;
output 	opcode_ex2;
output 	opcode_ex3;
output 	opcode_ex4;
input 	Equal131;
output 	memren_ex;
output 	memwen_ex;
output 	rdat1_mem1;
output 	pc_bran_mem1;
output 	rdat1_mem2;
output 	pc_bran_mem2;
output 	rdat1_mem3;
output 	pc_bran_mem3;
output 	rdat1_mem4;
output 	pc_bran_mem4;
output 	rdat1_mem5;
output 	pc_bran_mem5;
output 	rdat1_mem6;
output 	pc_bran_mem6;
output 	rdat1_mem7;
output 	pc_bran_mem7;
output 	rdat1_mem8;
output 	pc_bran_mem8;
output 	instr_mem6;
output 	rdat1_mem9;
output 	pc_bran_mem9;
output 	instr_mem7;
output 	rdat1_mem10;
output 	pc_bran_mem10;
output 	instr_mem8;
output 	rdat1_mem11;
output 	pc_bran_mem11;
output 	instr_mem9;
output 	rdat1_mem12;
output 	pc_bran_mem12;
output 	instr_mem10;
output 	rdat1_mem13;
output 	pc_bran_mem13;
output 	instr_mem11;
output 	rdat1_mem14;
output 	pc_bran_mem14;
output 	instr_mem12;
output 	rdat1_mem15;
output 	pc_bran_mem15;
output 	instr_mem13;
output 	rdat1_mem16;
output 	pc_bran_mem16;
output 	instr_mem14;
output 	rdat1_mem17;
output 	pc_bran_mem17;
output 	instr_mem15;
output 	rdat1_mem18;
output 	pc_bran_mem18;
output 	instr_mem16;
output 	rdat1_mem19;
output 	pc_bran_mem19;
input 	prifpc_mem_151;
output 	prifpc_mem_291;
output 	rdat1_mem20;
output 	pc_bran_mem20;
output 	prifpc_mem_281;
output 	rdat1_mem21;
output 	pc_bran_mem21;
output 	prifpc_mem_311;
output 	rdat1_mem22;
output 	pc_bran_mem22;
output 	prifpc_mem_301;
output 	rdat1_mem23;
output 	pc_bran_mem23;
output 	instr_mem17;
output 	rdat1_mem24;
output 	pc_bran_mem24;
output 	instr_mem18;
output 	rdat1_mem25;
output 	pc_bran_mem25;
output 	instr_mem19;
output 	rdat1_mem26;
output 	pc_bran_mem26;
output 	instr_mem20;
output 	rdat1_mem27;
output 	pc_bran_mem27;
output 	instr_mem21;
output 	rdat1_mem28;
output 	pc_bran_mem28;
output 	instr_mem22;
output 	rdat1_mem29;
output 	pc_bran_mem29;
output 	instr_mem23;
output 	rdat1_mem30;
output 	pc_bran_mem30;
output 	instr_mem24;
output 	rdat1_mem31;
output 	pc_bran_mem31;
output 	instr_mem25;
output 	dmemstore1;
output 	dmemstore2;
input 	Mux602;
output 	dmemstore3;
input 	Mux592;
output 	dmemstore4;
input 	Mux582;
output 	dmemstore5;
input 	Mux572;
output 	dmemstore6;
input 	Mux562;
output 	dmemstore7;
input 	Mux552;
output 	dmemstore8;
input 	Mux542;
output 	dmemstore9;
input 	Mux532;
output 	dmemstore10;
input 	Mux522;
output 	dmemstore11;
input 	Mux512;
output 	dmemstore12;
input 	Mux502;
output 	dmemstore13;
input 	Mux492;
output 	dmemstore14;
input 	Mux482;
output 	dmemstore15;
output 	dmemstore16;
output 	dmemstore17;
output 	dmemstore18;
output 	dmemstore19;
output 	dmemstore20;
output 	dmemstore21;
output 	dmemstore22;
output 	dmemstore23;
output 	dmemstore24;
output 	dmemstore25;
output 	dmemstore26;
output 	dmemstore27;
output 	dmemstore28;
output 	dmemstore29;
output 	dmemstore30;
output 	dmemstore31;
output 	halt_ex;
input 	prifhalt_wb;
input 	ifid_en;
output 	imemload_id;
output 	imemload_id1;
output 	imemload_id2;
output 	imemload_id3;
output 	imemload_id4;
output 	imemload_id5;
output 	imemload_id6;
output 	imemload_id7;
output 	imemload_id8;
output 	imemload_id9;
output 	imemload_id10;
output 	imemload_id11;
output 	imemload_id12;
output 	Regwen_ex;
output 	rd_ex;
output 	RegDest_ex;
output 	RegDest_ex1;
output 	rd_ex1;
output 	rd_ex2;
output 	rd_ex3;
output 	rd_ex4;
output 	imemload_id13;
output 	imemload_id14;
output 	imemload_id15;
output 	imemload_id16;
output 	imemload_id17;
output 	dataScr_mem;
output 	dataScr_mem1;
output 	prifpc_mem_110;
output 	imemload_id18;
output 	imemload_id19;
output 	imemload_id20;
output 	imemload_id21;
output 	imemload_id22;
output 	opcode_ex5;
output 	imemload_id23;
output 	prifpc_mem_01;
output 	prifpc_mem_32;
output 	imemload_id24;
output 	imemload_id25;
output 	prifpc_mem_210;
output 	prifpc_mem_41;
output 	imemload_id26;
output 	imemload_id27;
output 	prifpc_mem_51;
output 	prifpc_mem_152;
output 	imemload_id28;
output 	prifpc_mem_141;
output 	imemload_id29;
output 	prifpc_mem_131;
output 	imemload_id30;
output 	prifpc_mem_121;
output 	imemload_id31;
output 	prifpc_mem_111;
output 	prifpc_mem_101;
output 	prifpc_mem_91;
output 	prifpc_mem_61;
output 	prifpc_mem_271;
output 	prifpc_mem_231;
output 	prifpc_mem_181;
output 	prifpc_mem_241;
output 	prifpc_mem_161;
output 	prifpc_mem_191;
output 	prifpc_mem_171;
output 	prifpc_mem_211;
output 	prifpc_mem_201;
output 	prifpc_mem_261;
output 	prifpc_mem_81;
output 	prifpc_mem_71;
output 	prifpc_mem_221;
output 	prifpc_mem_251;
output 	instr_ex1;
output 	instr_ex2;
output 	instr_ex3;
output 	instr_ex4;
output 	instr_ex5;
output 	instr_ex6;
output 	PCScr_ex;
output 	pc_ex;
output 	PCScr_ex1;
output 	pc_ex1;
output 	pc_ex2;
output 	pc_ex3;
output 	pc_ex4;
output 	pc_ex5;
output 	pc_ex6;
output 	pc_ex7;
output 	pc_ex8;
output 	pc_ex9;
output 	instr_ex7;
output 	instr_ex8;
output 	pc_ex10;
output 	pc_ex11;
output 	instr_ex9;
output 	instr_ex10;
output 	pc_ex12;
output 	pc_ex13;
output 	instr_ex11;
output 	instr_ex12;
output 	pc_ex14;
output 	pc_ex15;
output 	instr_ex13;
output 	instr_ex14;
output 	pc_ex16;
output 	pc_ex17;
output 	pc_ex18;
output 	pc_ex19;
output 	pc_ex20;
output 	pc_ex21;
output 	pc_ex22;
output 	pc_ex23;
output 	instr_ex15;
output 	instr_ex16;
output 	instr_ex17;
output 	pc_ex24;
output 	pc_ex25;
output 	pc_ex26;
output 	pc_ex27;
output 	pc_ex28;
output 	pc_ex29;
output 	pc_ex30;
output 	pc_ex31;
output 	instr_ex18;
output 	instr_ex19;
output 	instr_ex20;
output 	instr_ex21;
output 	instr_ex22;
output 	instr_ex23;
output 	instr_ex24;
output 	instr_ex25;
output 	halt_wb;
output 	dataScr_ex1;
output 	pc_id;
output 	pc_id1;
output 	pc_id2;
output 	pc_id3;
output 	pc_id4;
output 	pc_id5;
output 	pc_id6;
output 	pc_id7;
output 	pc_id8;
output 	pc_id9;
output 	pc_id10;
output 	pc_id11;
output 	pc_id12;
output 	pc_id13;
output 	pc_id14;
output 	pc_id15;
output 	pc_id16;
output 	pc_id17;
output 	pc_id18;
output 	pc_id19;
output 	pc_id20;
output 	pc_id21;
output 	pc_id22;
output 	pc_id23;
output 	pc_id24;
output 	pc_id25;
output 	pc_id26;
output 	pc_id27;
output 	pc_id28;
output 	pc_id29;
output 	pc_id30;
output 	pc_id31;
output 	dataScr_ex2;
output 	ALUScr_ex3;
output 	zero_flag_mem;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \zero_flag_mem~3_combout ;
wire \zero_flag_mem~4_combout ;
wire \zero_flag_mem~5_combout ;
wire \zero_flag_mem~8_combout ;
wire \ALUScr_ex~10_combout ;
wire \ALUScr_ex~14_combout ;
wire \ALUScr_ex~9_combout ;
wire \regwrite_mem~0_combout ;
wire \regwrite_mem~2_combout ;
wire \regwrite_mem~4_combout ;
wire \regwrite_mem~6_combout ;
wire \regwrite_mem~8_combout ;
wire \rdat2_ex~0_combout ;
wire \rdat1_ex~0_combout ;
wire \rdat2_ex~2_combout ;
wire \rdat1_ex~2_combout ;
wire \rdat2_ex~4_combout ;
wire \rdat2_ex~6_combout ;
wire \rdat2_ex~8_combout ;
wire \rdat2_ex~10_combout ;
wire \rdat2_ex~12_combout ;
wire \rdat2_ex~14_combout ;
wire \rdat2_ex~16_combout ;
wire \rdat2_ex~18_combout ;
wire \rdat2_ex~20_combout ;
wire \rdat2_ex~22_combout ;
wire \rdat2_ex~24_combout ;
wire \rdat2_ex~26_combout ;
wire \rdat2_ex~28_combout ;
wire \rdat2_ex~30_combout ;
wire \rdat2_ex~32_combout ;
wire \rdat2_ex~34_combout ;
wire \rdat2_ex~36_combout ;
wire \rdat2_ex~38_combout ;
wire \rdat2_ex~40_combout ;
wire \rdat2_ex~42_combout ;
wire \rdat2_ex~44_combout ;
wire \rdat2_ex~46_combout ;
wire \rdat2_ex~48_combout ;
wire \rdat2_ex~50_combout ;
wire \rdat2_ex~52_combout ;
wire \rdat2_ex~54_combout ;
wire \rdat2_ex~56_combout ;
wire \rdat2_ex~58_combout ;
wire \rdat2_ex~60_combout ;
wire \rdat2_ex~62_combout ;
wire \ALUOP_ex~1_combout ;
wire \rdat1_ex~4_combout ;
wire \rdat1_ex~6_combout ;
wire \rdat1_ex~8_combout ;
wire \rdat1_ex~10_combout ;
wire \rdat1_ex~12_combout ;
wire \rdat1_ex~14_combout ;
wire \rdat1_ex~16_combout ;
wire \rdat1_ex~18_combout ;
wire \rdat1_ex~20_combout ;
wire \rdat1_ex~22_combout ;
wire \rdat1_ex~24_combout ;
wire \rdat1_ex~26_combout ;
wire \rdat1_ex~28_combout ;
wire \rdat1_ex~30_combout ;
wire \rdat1_ex~32_combout ;
wire \rdat1_ex~34_combout ;
wire \rdat1_ex~36_combout ;
wire \rdat1_ex~38_combout ;
wire \rdat1_ex~40_combout ;
wire \rdat1_ex~42_combout ;
wire \rdat1_ex~44_combout ;
wire \rdat1_ex~46_combout ;
wire \rdat1_ex~48_combout ;
wire \rdat1_ex~50_combout ;
wire \rdat1_ex~52_combout ;
wire \rdat1_ex~54_combout ;
wire \rdat1_ex~56_combout ;
wire \rdat1_ex~58_combout ;
wire \rdat1_ex~60_combout ;
wire \rdat1_ex~62_combout ;
wire \PCScr_ex~2_combout ;
wire \PCScr_ex~5_combout ;
wire \ALUScr_ex~5_combout ;
wire \ALUScr_ex~6_combout ;
wire \zero_flag_mem~0_combout ;
wire \zero_flag_mem~6_combout ;
wire \zero_flag_mem~9_combout ;
wire \zero_flag_mem~7_combout ;
wire \zero_flag_mem~10_combout ;
wire \zero_flag_mem~11_combout ;
wire \zero_flag_mem~12_combout ;
wire \zero_flag_mem~1_combout ;
wire \zero_flag_mem~2_combout ;


// Location: LCCOMB_X60_Y25_N20
cycloneive_lcell_comb \zero_flag_mem~3 (
// Equation(s):
// \zero_flag_mem~3_combout  = (!aluifportOut_6 & (!aluifportOut_53 & ((!aluifportOut_51) # (!aluifportOut_5))))

	.dataa(aluifportOut_6),
	.datab(aluifportOut_5),
	.datac(aluifportOut_51),
	.datad(aluifportOut_53),
	.cin(gnd),
	.combout(\zero_flag_mem~3_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~3 .lut_mask = 16'h0015;
defparam \zero_flag_mem~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N6
cycloneive_lcell_comb \zero_flag_mem~4 (
// Equation(s):
// \zero_flag_mem~4_combout  = (!aluifportOut_26 & (!aluifportOut_24 & (!aluifportOut_25 & !aluifportOut_27)))

	.dataa(aluifportOut_26),
	.datab(aluifportOut_24),
	.datac(aluifportOut_25),
	.datad(aluifportOut_27),
	.cin(gnd),
	.combout(\zero_flag_mem~4_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~4 .lut_mask = 16'h0001;
defparam \zero_flag_mem~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N22
cycloneive_lcell_comb \zero_flag_mem~5 (
// Equation(s):
// \zero_flag_mem~5_combout  = (!aluifportOut_4 & (\zero_flag_mem~4_combout  & (!aluifportOut_7 & \zero_flag_mem~3_combout )))

	.dataa(aluifportOut_4),
	.datab(\zero_flag_mem~4_combout ),
	.datac(aluifportOut_7),
	.datad(\zero_flag_mem~3_combout ),
	.cin(gnd),
	.combout(\zero_flag_mem~5_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~5 .lut_mask = 16'h0400;
defparam \zero_flag_mem~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N26
cycloneive_lcell_comb \zero_flag_mem~8 (
// Equation(s):
// \zero_flag_mem~8_combout  = ((!aluifportOut_8 & (!aluifportOut_23 & !aluifportOut_12))) # (!\prif.ALUOP_ex [3])

	.dataa(prifALUOP_ex_3),
	.datab(aluifportOut_8),
	.datac(aluifportOut_23),
	.datad(aluifportOut_12),
	.cin(gnd),
	.combout(\zero_flag_mem~8_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~8 .lut_mask = 16'h5557;
defparam \zero_flag_mem~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N24
cycloneive_lcell_comb \dmemaddr~0 (
// Equation(s):
// dmemaddr = (exmem_en & ((aluifportOut_1))) # (!exmem_en & (prifdmemaddr_1))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemaddr_1),
	.datad(aluifportOut_1),
	.cin(gnd),
	.combout(dmemaddr),
	.cout());
// synopsys translate_off
defparam \dmemaddr~0 .lut_mask = 16'hFA50;
defparam \dmemaddr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N28
cycloneive_lcell_comb \dmemren~0 (
// Equation(s):
// dmemren = (prifdmemren) # ((\prif.memren_ex~q  & exmem_en))

	.dataa(prifmemren_ex),
	.datab(gnd),
	.datac(prifdmemren),
	.datad(exmem_en),
	.cin(gnd),
	.combout(dmemren),
	.cout());
// synopsys translate_off
defparam \dmemren~0 .lut_mask = 16'hFAF0;
defparam \dmemren~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N14
cycloneive_lcell_comb \dmemwen~0 (
// Equation(s):
// dmemwen = (prifdmemwen) # ((\prif.memwen_ex~q  & exmem_en))

	.dataa(prifmemwen_ex),
	.datab(gnd),
	.datac(prifdmemwen),
	.datad(exmem_en),
	.cin(gnd),
	.combout(dmemwen),
	.cout());
// synopsys translate_off
defparam \dmemwen~0 .lut_mask = 16'hFAF0;
defparam \dmemwen~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N4
cycloneive_lcell_comb \dmemaddr~1 (
// Equation(s):
// dmemaddr1 = (exmem_en & (aluifportOut_0)) # (!exmem_en & ((prifdmemaddr_0)))

	.dataa(gnd),
	.datab(aluifportOut_0),
	.datac(prifdmemaddr_0),
	.datad(exmem_en),
	.cin(gnd),
	.combout(dmemaddr1),
	.cout());
// synopsys translate_off
defparam \dmemaddr~1 .lut_mask = 16'hCCF0;
defparam \dmemaddr~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N30
cycloneive_lcell_comb \dmemaddr~2 (
// Equation(s):
// dmemaddr2 = (exmem_en & ((aluifportOut_32))) # (!exmem_en & (prifdmemaddr_3))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemaddr_3),
	.datad(aluifportOut_32),
	.cin(gnd),
	.combout(dmemaddr2),
	.cout());
// synopsys translate_off
defparam \dmemaddr~2 .lut_mask = 16'hFA50;
defparam \dmemaddr~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N0
cycloneive_lcell_comb \dmemaddr~3 (
// Equation(s):
// dmemaddr3 = (exmem_en & (aluifportOut_21)) # (!exmem_en & ((prifdmemaddr_2)))

	.dataa(gnd),
	.datab(aluifportOut_21),
	.datac(prifdmemaddr_2),
	.datad(exmem_en),
	.cin(gnd),
	.combout(dmemaddr3),
	.cout());
// synopsys translate_off
defparam \dmemaddr~3 .lut_mask = 16'hCCF0;
defparam \dmemaddr~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N16
cycloneive_lcell_comb \dmemaddr~4 (
// Equation(s):
// dmemaddr4 = (exmem_en & ((aluifportOut_52))) # (!exmem_en & (prifdmemaddr_5))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemaddr_5),
	.datad(aluifportOut_52),
	.cin(gnd),
	.combout(dmemaddr4),
	.cout());
// synopsys translate_off
defparam \dmemaddr~4 .lut_mask = 16'hFA50;
defparam \dmemaddr~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N18
cycloneive_lcell_comb \dmemaddr~5 (
// Equation(s):
// dmemaddr5 = (exmem_en & (aluifportOut_4)) # (!exmem_en & ((prifdmemaddr_4)))

	.dataa(gnd),
	.datab(aluifportOut_4),
	.datac(prifdmemaddr_4),
	.datad(exmem_en),
	.cin(gnd),
	.combout(dmemaddr5),
	.cout());
// synopsys translate_off
defparam \dmemaddr~5 .lut_mask = 16'hCCF0;
defparam \dmemaddr~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N4
cycloneive_lcell_comb \dmemaddr~6 (
// Equation(s):
// dmemaddr6 = (exmem_en & ((aluifportOut_7))) # (!exmem_en & (prifdmemaddr_7))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemaddr_7),
	.datad(aluifportOut_7),
	.cin(gnd),
	.combout(dmemaddr6),
	.cout());
// synopsys translate_off
defparam \dmemaddr~6 .lut_mask = 16'hFA50;
defparam \dmemaddr~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N14
cycloneive_lcell_comb \dmemaddr~7 (
// Equation(s):
// dmemaddr7 = (exmem_en & ((aluifportOut_6))) # (!exmem_en & (prifdmemaddr_6))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemaddr_6),
	.datad(aluifportOut_6),
	.cin(gnd),
	.combout(dmemaddr7),
	.cout());
// synopsys translate_off
defparam \dmemaddr~7 .lut_mask = 16'hFA50;
defparam \dmemaddr~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N8
cycloneive_lcell_comb \dmemaddr~8 (
// Equation(s):
// dmemaddr8 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_9)))) # (!exmem_en & (((prifdmemaddr_9))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_9),
	.datad(aluifportOut_9),
	.cin(gnd),
	.combout(dmemaddr8),
	.cout());
// synopsys translate_off
defparam \dmemaddr~8 .lut_mask = 16'hD850;
defparam \dmemaddr~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N22
cycloneive_lcell_comb \dmemaddr~9 (
// Equation(s):
// dmemaddr9 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_8)))) # (!exmem_en & (((prifdmemaddr_8))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_8),
	.datad(aluifportOut_8),
	.cin(gnd),
	.combout(dmemaddr9),
	.cout());
// synopsys translate_off
defparam \dmemaddr~9 .lut_mask = 16'hD850;
defparam \dmemaddr~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N22
cycloneive_lcell_comb \dmemaddr~10 (
// Equation(s):
// dmemaddr10 = (exmem_en & (\prif.ALUOP_ex [3] & (aluifportOut_11))) # (!exmem_en & (((prifdmemaddr_11))))

	.dataa(prifALUOP_ex_3),
	.datab(aluifportOut_11),
	.datac(prifdmemaddr_11),
	.datad(exmem_en),
	.cin(gnd),
	.combout(dmemaddr10),
	.cout());
// synopsys translate_off
defparam \dmemaddr~10 .lut_mask = 16'h88F0;
defparam \dmemaddr~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N16
cycloneive_lcell_comb \dmemaddr~11 (
// Equation(s):
// dmemaddr11 = (exmem_en & (\prif.ALUOP_ex [3] & (aluifportOut_10))) # (!exmem_en & (((prifdmemaddr_10))))

	.dataa(prifALUOP_ex_3),
	.datab(aluifportOut_10),
	.datac(prifdmemaddr_10),
	.datad(exmem_en),
	.cin(gnd),
	.combout(dmemaddr11),
	.cout());
// synopsys translate_off
defparam \dmemaddr~11 .lut_mask = 16'h88F0;
defparam \dmemaddr~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N12
cycloneive_lcell_comb \dmemaddr~12 (
// Equation(s):
// dmemaddr12 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_13)))) # (!exmem_en & (((prifdmemaddr_13))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_13),
	.datad(aluifportOut_13),
	.cin(gnd),
	.combout(dmemaddr12),
	.cout());
// synopsys translate_off
defparam \dmemaddr~12 .lut_mask = 16'hD850;
defparam \dmemaddr~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N30
cycloneive_lcell_comb \dmemaddr~13 (
// Equation(s):
// dmemaddr13 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_12)))) # (!exmem_en & (((prifdmemaddr_12))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_12),
	.datad(aluifportOut_12),
	.cin(gnd),
	.combout(dmemaddr13),
	.cout());
// synopsys translate_off
defparam \dmemaddr~13 .lut_mask = 16'hD850;
defparam \dmemaddr~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N8
cycloneive_lcell_comb \dmemaddr~14 (
// Equation(s):
// dmemaddr14 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_15)))) # (!exmem_en & (((prifdmemaddr_15))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_15),
	.datad(aluifportOut_15),
	.cin(gnd),
	.combout(dmemaddr14),
	.cout());
// synopsys translate_off
defparam \dmemaddr~14 .lut_mask = 16'hD850;
defparam \dmemaddr~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N8
cycloneive_lcell_comb \dmemaddr~15 (
// Equation(s):
// dmemaddr15 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_14)))) # (!exmem_en & (((prifdmemaddr_14))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_14),
	.datad(aluifportOut_14),
	.cin(gnd),
	.combout(dmemaddr15),
	.cout());
// synopsys translate_off
defparam \dmemaddr~15 .lut_mask = 16'hD850;
defparam \dmemaddr~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N4
cycloneive_lcell_comb \dmemaddr~16 (
// Equation(s):
// dmemaddr16 = (exmem_en & (aluifportOut_23 & ((\prif.ALUOP_ex [3])))) # (!exmem_en & (((prifdmemaddr_23))))

	.dataa(aluifportOut_23),
	.datab(exmem_en),
	.datac(prifdmemaddr_23),
	.datad(prifALUOP_ex_3),
	.cin(gnd),
	.combout(dmemaddr16),
	.cout());
// synopsys translate_off
defparam \dmemaddr~16 .lut_mask = 16'hB830;
defparam \dmemaddr~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N14
cycloneive_lcell_comb \dmemaddr~17 (
// Equation(s):
// dmemaddr17 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_22)))) # (!exmem_en & (((prifdmemaddr_22))))

	.dataa(prifALUOP_ex_3),
	.datab(exmem_en),
	.datac(prifdmemaddr_22),
	.datad(aluifportOut_22),
	.cin(gnd),
	.combout(dmemaddr17),
	.cout());
// synopsys translate_off
defparam \dmemaddr~17 .lut_mask = 16'hB830;
defparam \dmemaddr~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N28
cycloneive_lcell_comb \dmemaddr~18 (
// Equation(s):
// dmemaddr18 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_211)))) # (!exmem_en & (((prifdmemaddr_21))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_21),
	.datad(aluifportOut_211),
	.cin(gnd),
	.combout(dmemaddr18),
	.cout());
// synopsys translate_off
defparam \dmemaddr~18 .lut_mask = 16'hD850;
defparam \dmemaddr~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N8
cycloneive_lcell_comb \dmemaddr~19 (
// Equation(s):
// dmemaddr19 = (exmem_en & ((aluifportOut_29))) # (!exmem_en & (prifdmemaddr_29))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemaddr_29),
	.datad(aluifportOut_29),
	.cin(gnd),
	.combout(dmemaddr19),
	.cout());
// synopsys translate_off
defparam \dmemaddr~19 .lut_mask = 16'hFA50;
defparam \dmemaddr~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N26
cycloneive_lcell_comb \dmemaddr~20 (
// Equation(s):
// dmemaddr20 = (exmem_en & ((aluifportOut_28))) # (!exmem_en & (prifdmemaddr_28))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemaddr_28),
	.datad(aluifportOut_28),
	.cin(gnd),
	.combout(dmemaddr20),
	.cout());
// synopsys translate_off
defparam \dmemaddr~20 .lut_mask = 16'hFA50;
defparam \dmemaddr~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N8
cycloneive_lcell_comb \dmemaddr~21 (
// Equation(s):
// dmemaddr21 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifneg_flag)))) # (!exmem_en & (((prifdmemaddr_31))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_31),
	.datad(aluifneg_flag),
	.cin(gnd),
	.combout(dmemaddr21),
	.cout());
// synopsys translate_off
defparam \dmemaddr~21 .lut_mask = 16'hD850;
defparam \dmemaddr~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N0
cycloneive_lcell_comb \dmemaddr~22 (
// Equation(s):
// dmemaddr22 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_30)))) # (!exmem_en & (((prifdmemaddr_30))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_30),
	.datad(aluifportOut_30),
	.cin(gnd),
	.combout(dmemaddr22),
	.cout());
// synopsys translate_off
defparam \dmemaddr~22 .lut_mask = 16'hD850;
defparam \dmemaddr~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N0
cycloneive_lcell_comb \dmemaddr~23 (
// Equation(s):
// dmemaddr23 = (exmem_en & (aluifportOut_20 & ((\prif.ALUOP_ex [3])))) # (!exmem_en & (((prifdmemaddr_20))))

	.dataa(aluifportOut_20),
	.datab(exmem_en),
	.datac(prifdmemaddr_20),
	.datad(prifALUOP_ex_3),
	.cin(gnd),
	.combout(dmemaddr23),
	.cout());
// synopsys translate_off
defparam \dmemaddr~23 .lut_mask = 16'hB830;
defparam \dmemaddr~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N10
cycloneive_lcell_comb \dmemaddr~24 (
// Equation(s):
// dmemaddr24 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_17)))) # (!exmem_en & (((prifdmemaddr_17))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_17),
	.datad(aluifportOut_17),
	.cin(gnd),
	.combout(dmemaddr24),
	.cout());
// synopsys translate_off
defparam \dmemaddr~24 .lut_mask = 16'hD850;
defparam \dmemaddr~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N12
cycloneive_lcell_comb \dmemaddr~25 (
// Equation(s):
// dmemaddr25 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_16)))) # (!exmem_en & (((prifdmemaddr_16))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_16),
	.datad(aluifportOut_16),
	.cin(gnd),
	.combout(dmemaddr25),
	.cout());
// synopsys translate_off
defparam \dmemaddr~25 .lut_mask = 16'hD850;
defparam \dmemaddr~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N0
cycloneive_lcell_comb \dmemaddr~26 (
// Equation(s):
// dmemaddr26 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_19)))) # (!exmem_en & (((prifdmemaddr_19))))

	.dataa(exmem_en),
	.datab(prifALUOP_ex_3),
	.datac(prifdmemaddr_19),
	.datad(aluifportOut_19),
	.cin(gnd),
	.combout(dmemaddr26),
	.cout());
// synopsys translate_off
defparam \dmemaddr~26 .lut_mask = 16'hD850;
defparam \dmemaddr~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y25_N4
cycloneive_lcell_comb \dmemaddr~27 (
// Equation(s):
// dmemaddr27 = (exmem_en & (\prif.ALUOP_ex [3] & ((aluifportOut_18)))) # (!exmem_en & (((prifdmemaddr_18))))

	.dataa(prifALUOP_ex_3),
	.datab(exmem_en),
	.datac(prifdmemaddr_18),
	.datad(aluifportOut_18),
	.cin(gnd),
	.combout(dmemaddr27),
	.cout());
// synopsys translate_off
defparam \dmemaddr~27 .lut_mask = 16'hB830;
defparam \dmemaddr~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N16
cycloneive_lcell_comb \dmemaddr~28 (
// Equation(s):
// dmemaddr28 = (exmem_en & ((aluifportOut_25))) # (!exmem_en & (prifdmemaddr_25))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemaddr_25),
	.datad(aluifportOut_25),
	.cin(gnd),
	.combout(dmemaddr28),
	.cout());
// synopsys translate_off
defparam \dmemaddr~28 .lut_mask = 16'hFA50;
defparam \dmemaddr~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N12
cycloneive_lcell_comb \dmemaddr~29 (
// Equation(s):
// dmemaddr29 = (exmem_en & ((aluifportOut_24))) # (!exmem_en & (prifdmemaddr_24))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemaddr_24),
	.datad(aluifportOut_24),
	.cin(gnd),
	.combout(dmemaddr29),
	.cout());
// synopsys translate_off
defparam \dmemaddr~29 .lut_mask = 16'hFA50;
defparam \dmemaddr~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N28
cycloneive_lcell_comb \dmemaddr~30 (
// Equation(s):
// dmemaddr30 = (exmem_en & ((aluifportOut_27))) # (!exmem_en & (prifdmemaddr_27))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemaddr_27),
	.datad(aluifportOut_27),
	.cin(gnd),
	.combout(dmemaddr30),
	.cout());
// synopsys translate_off
defparam \dmemaddr~30 .lut_mask = 16'hFC30;
defparam \dmemaddr~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N12
cycloneive_lcell_comb \dmemaddr~31 (
// Equation(s):
// dmemaddr31 = (exmem_en & ((aluifportOut_26))) # (!exmem_en & (prifdmemaddr_26))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemaddr_26),
	.datad(aluifportOut_26),
	.cin(gnd),
	.combout(dmemaddr31),
	.cout());
// synopsys translate_off
defparam \dmemaddr~31 .lut_mask = 16'hFC30;
defparam \dmemaddr~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N24
cycloneive_lcell_comb \halt_mem~0 (
// Equation(s):
// halt_mem = (exmem_en & ((\prif.halt_ex~q ))) # (!exmem_en & (\prif.halt_mem~q ))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifhalt_mem),
	.datad(prifhalt_ex),
	.cin(gnd),
	.combout(halt_mem),
	.cout());
// synopsys translate_off
defparam \halt_mem~0 .lut_mask = 16'hFC30;
defparam \halt_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N10
cycloneive_lcell_comb \dmemstore~0 (
// Equation(s):
// dmemstore = (exmem_en & ((\Mux63~1_combout ) # ((\Mux63~0_combout )))) # (!exmem_en & (((prifdmemstore_0))))

	.dataa(Mux631),
	.datab(exmem_en),
	.datac(prifdmemstore_0),
	.datad(Mux63),
	.cin(gnd),
	.combout(dmemstore),
	.cout());
// synopsys translate_off
defparam \dmemstore~0 .lut_mask = 16'hFCB8;
defparam \dmemstore~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N0
cycloneive_lcell_comb \dataScr_ex~2 (
// Equation(s):
// dataScr_ex = (!Equal13 & (((!\prif.imemload_id [26]) # (!\prif.imemload_id [27])) # (!Equal20)))

	.dataa(Equal20),
	.datab(prifimemload_id_27),
	.datac(prifimemload_id_26),
	.datad(Equal13),
	.cin(gnd),
	.combout(dataScr_ex),
	.cout());
// synopsys translate_off
defparam \dataScr_ex~2 .lut_mask = 16'h007F;
defparam \dataScr_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N14
cycloneive_lcell_comb \ALUOP_ex~0 (
// Equation(s):
// ALUOP_ex = (!flush_idex & ((ccifiwait_0 & (\prif.ALUOP_ex [3])) # (!ccifiwait_0 & ((!Selector0)))))

	.dataa(ccifiwait_0),
	.datab(flush_idex),
	.datac(prifALUOP_ex_3),
	.datad(Selector0),
	.cin(gnd),
	.combout(ALUOP_ex),
	.cout());
// synopsys translate_off
defparam \ALUOP_ex~0 .lut_mask = 16'h2031;
defparam \ALUOP_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N28
cycloneive_lcell_comb \imm_ex~0 (
// Equation(s):
// imm_ex = (ccifiwait_0 & (\prif.imm_ex [1])) # (!ccifiwait_0 & ((\prif.imemload_id [1])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifimm_ex_1),
	.datad(prifimemload_id_1),
	.cin(gnd),
	.combout(imm_ex),
	.cout());
// synopsys translate_off
defparam \imm_ex~0 .lut_mask = 16'hF5A0;
defparam \imm_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N4
cycloneive_lcell_comb \ALUScr_ex~11 (
// Equation(s):
// ALUScr_ex = (ccifiwait_0 & ((\prif.ALUScr_ex [1]))) # (!ccifiwait_0 & (\ALUScr_ex~14_combout ))

	.dataa(ccifiwait_0),
	.datab(\ALUScr_ex~14_combout ),
	.datac(prifALUScr_ex_1),
	.datad(gnd),
	.cin(gnd),
	.combout(ALUScr_ex),
	.cout());
// synopsys translate_off
defparam \ALUScr_ex~11 .lut_mask = 16'hE4E4;
defparam \ALUScr_ex~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N30
cycloneive_lcell_comb \shamt_ex~0 (
// Equation(s):
// shamt_ex = (ccifiwait_0 & ((\prif.shamt_ex [1]))) # (!ccifiwait_0 & (\prif.imemload_id [7]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_7),
	.datac(prifshamt_ex_1),
	.datad(gnd),
	.cin(gnd),
	.combout(shamt_ex),
	.cout());
// synopsys translate_off
defparam \shamt_ex~0 .lut_mask = 16'hE4E4;
defparam \shamt_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N20
cycloneive_lcell_comb \ALUScr_ex~12 (
// Equation(s):
// ALUScr_ex1 = (ccifiwait_0 & (\prif.ALUScr_ex [0])) # (!ccifiwait_0 & (((ALUScr_ex3 & \ALUScr_ex~9_combout ))))

	.dataa(prifALUScr_ex_0),
	.datab(ALUScr_ex3),
	.datac(\ALUScr_ex~9_combout ),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(ALUScr_ex1),
	.cout());
// synopsys translate_off
defparam \ALUScr_ex~12 .lut_mask = 16'hAAC0;
defparam \ALUScr_ex~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N12
cycloneive_lcell_comb \Regwen_mem~0 (
// Equation(s):
// Regwen_mem = (exmem_en & (\prif.Regwen_ex~q )) # (!exmem_en & ((\prif.Regwen_mem~q )))

	.dataa(gnd),
	.datab(prifRegwen_ex),
	.datac(prifRegwen_mem),
	.datad(exmem_en),
	.cin(gnd),
	.combout(Regwen_mem),
	.cout());
// synopsys translate_off
defparam \Regwen_mem~0 .lut_mask = 16'hCCF0;
defparam \Regwen_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N10
cycloneive_lcell_comb \regwrite_mem~1 (
// Equation(s):
// regwrite_mem = (exmem_en & (\regwrite_mem~0_combout )) # (!exmem_en & ((\prif.regwrite_mem [4])))

	.dataa(\regwrite_mem~0_combout ),
	.datab(exmem_en),
	.datac(prifregwrite_mem_4),
	.datad(gnd),
	.cin(gnd),
	.combout(regwrite_mem),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~1 .lut_mask = 16'hB8B8;
defparam \regwrite_mem~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N4
cycloneive_lcell_comb \regwrite_mem~3 (
// Equation(s):
// regwrite_mem1 = (exmem_en & ((\regwrite_mem~2_combout ))) # (!exmem_en & (\prif.regwrite_mem [0]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifregwrite_mem_0),
	.datad(\regwrite_mem~2_combout ),
	.cin(gnd),
	.combout(regwrite_mem1),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~3 .lut_mask = 16'hFC30;
defparam \regwrite_mem~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N26
cycloneive_lcell_comb \regwrite_mem~5 (
// Equation(s):
// regwrite_mem2 = (exmem_en & ((\regwrite_mem~4_combout ))) # (!exmem_en & (\prif.regwrite_mem [1]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifregwrite_mem_1),
	.datad(\regwrite_mem~4_combout ),
	.cin(gnd),
	.combout(regwrite_mem2),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~5 .lut_mask = 16'hFC30;
defparam \regwrite_mem~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N0
cycloneive_lcell_comb \regwrite_mem~7 (
// Equation(s):
// regwrite_mem3 = (exmem_en & ((\regwrite_mem~6_combout ))) # (!exmem_en & (\prif.regwrite_mem [2]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifregwrite_mem_2),
	.datad(\regwrite_mem~6_combout ),
	.cin(gnd),
	.combout(regwrite_mem3),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~7 .lut_mask = 16'hFC30;
defparam \regwrite_mem~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N22
cycloneive_lcell_comb \regwrite_mem~9 (
// Equation(s):
// regwrite_mem4 = (exmem_en & ((\regwrite_mem~8_combout ))) # (!exmem_en & (\prif.regwrite_mem [3]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifregwrite_mem_3),
	.datad(\regwrite_mem~8_combout ),
	.cin(gnd),
	.combout(regwrite_mem4),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~9 .lut_mask = 16'hFC30;
defparam \regwrite_mem~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N24
cycloneive_lcell_comb \rt_ex~0 (
// Equation(s):
// rt_ex = (ccifiwait_0 & (\prif.rt_ex [1])) # (!ccifiwait_0 & ((\prif.imemload_id [17])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrt_ex_1),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(rt_ex),
	.cout());
// synopsys translate_off
defparam \rt_ex~0 .lut_mask = 16'hF3C0;
defparam \rt_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N2
cycloneive_lcell_comb \rt_ex~1 (
// Equation(s):
// rt_ex1 = (ccifiwait_0 & (\prif.rt_ex [0])) # (!ccifiwait_0 & ((\prif.imemload_id [16])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrt_ex_0),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(rt_ex1),
	.cout());
// synopsys translate_off
defparam \rt_ex~1 .lut_mask = 16'hF3C0;
defparam \rt_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N4
cycloneive_lcell_comb \rt_ex~2 (
// Equation(s):
// rt_ex2 = (ccifiwait_0 & (\prif.rt_ex [3])) # (!ccifiwait_0 & ((\prif.imemload_id [19])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrt_ex_3),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(rt_ex2),
	.cout());
// synopsys translate_off
defparam \rt_ex~2 .lut_mask = 16'hF3C0;
defparam \rt_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N10
cycloneive_lcell_comb \rt_ex~3 (
// Equation(s):
// rt_ex3 = (ccifiwait_0 & (\prif.rt_ex [2])) # (!ccifiwait_0 & ((\prif.imemload_id [18])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrt_ex_2),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(rt_ex3),
	.cout());
// synopsys translate_off
defparam \rt_ex~3 .lut_mask = 16'hF3C0;
defparam \rt_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y27_N8
cycloneive_lcell_comb \rt_ex~4 (
// Equation(s):
// rt_ex4 = (ccifiwait_0 & ((\prif.rt_ex [4]))) # (!ccifiwait_0 & (\prif.imemload_id [20]))

	.dataa(prifimemload_id_20),
	.datab(ccifiwait_0),
	.datac(prifrt_ex_4),
	.datad(gnd),
	.cin(gnd),
	.combout(rt_ex4),
	.cout());
// synopsys translate_off
defparam \rt_ex~4 .lut_mask = 16'hE2E2;
defparam \rt_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N2
cycloneive_lcell_comb \Regwen_wb~0 (
// Equation(s):
// Regwen_wb = (always1 & (\prif.Regwen_mem~q )) # (!always1 & ((\prif.Regwen_wb~q )))

	.dataa(prifRegwen_mem),
	.datab(gnd),
	.datac(prifRegwen_wb),
	.datad(always1),
	.cin(gnd),
	.combout(Regwen_wb),
	.cout());
// synopsys translate_off
defparam \Regwen_wb~0 .lut_mask = 16'hAAF0;
defparam \Regwen_wb~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N28
cycloneive_lcell_comb \regwrite_wb~0 (
// Equation(s):
// regwrite_wb = (always1 & ((\prif.regwrite_mem [2]))) # (!always1 & (\prif.regwrite_wb [2]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifregwrite_wb_2),
	.datad(prifregwrite_mem_2),
	.cin(gnd),
	.combout(regwrite_wb),
	.cout());
// synopsys translate_off
defparam \regwrite_wb~0 .lut_mask = 16'hFA50;
defparam \regwrite_wb~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N18
cycloneive_lcell_comb \regwrite_wb~1 (
// Equation(s):
// regwrite_wb1 = (always1 & (\prif.regwrite_mem [0])) # (!always1 & ((\prif.regwrite_wb [0])))

	.dataa(gnd),
	.datab(prifregwrite_mem_0),
	.datac(prifregwrite_wb_0),
	.datad(always1),
	.cin(gnd),
	.combout(regwrite_wb1),
	.cout());
// synopsys translate_off
defparam \regwrite_wb~1 .lut_mask = 16'hCCF0;
defparam \regwrite_wb~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N28
cycloneive_lcell_comb \regwrite_wb~2 (
// Equation(s):
// regwrite_wb2 = (always1 & (\prif.regwrite_mem [1])) # (!always1 & ((\prif.regwrite_wb [1])))

	.dataa(prifregwrite_mem_1),
	.datab(gnd),
	.datac(prifregwrite_wb_1),
	.datad(always1),
	.cin(gnd),
	.combout(regwrite_wb2),
	.cout());
// synopsys translate_off
defparam \regwrite_wb~2 .lut_mask = 16'hAAF0;
defparam \regwrite_wb~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N24
cycloneive_lcell_comb \regwrite_wb~3 (
// Equation(s):
// regwrite_wb3 = (always1 & (\prif.regwrite_mem [4])) # (!always1 & ((\prif.regwrite_wb [4])))

	.dataa(prifregwrite_mem_4),
	.datab(gnd),
	.datac(prifregwrite_wb_4),
	.datad(always1),
	.cin(gnd),
	.combout(regwrite_wb3),
	.cout());
// synopsys translate_off
defparam \regwrite_wb~3 .lut_mask = 16'hAAF0;
defparam \regwrite_wb~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N14
cycloneive_lcell_comb \regwrite_wb~4 (
// Equation(s):
// regwrite_wb4 = (always1 & (\prif.regwrite_mem [3])) # (!always1 & ((\prif.regwrite_wb [3])))

	.dataa(prifregwrite_mem_3),
	.datab(gnd),
	.datac(prifregwrite_wb_3),
	.datad(always1),
	.cin(gnd),
	.combout(regwrite_wb4),
	.cout());
// synopsys translate_off
defparam \regwrite_wb~4 .lut_mask = 16'hAAF0;
defparam \regwrite_wb~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N22
cycloneive_lcell_comb \dmemload_wb~0 (
// Equation(s):
// dmemload_wb = (always1 & (ramiframload_1)) # (!always1 & ((\prif.dmemload_wb [1])))

	.dataa(always1),
	.datab(ramiframload_1),
	.datac(prifdmemload_wb_1),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemload_wb),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~0 .lut_mask = 16'hD8D8;
defparam \dmemload_wb~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N20
cycloneive_lcell_comb \dmemaddr_wb~0 (
// Equation(s):
// dmemaddr_wb = (always1 & ((prifdmemaddr_1))) # (!always1 & (\prif.dmemaddr_wb [1]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_1),
	.datad(prifdmemaddr_1),
	.cin(gnd),
	.combout(dmemaddr_wb),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~0 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N6
cycloneive_lcell_comb \dataScr_wb~0 (
// Equation(s):
// dataScr_wb = (always1 & (\prif.dataScr_mem [0])) # (!always1 & ((\prif.dataScr_wb [0])))

	.dataa(prifdataScr_mem_0),
	.datab(gnd),
	.datac(prifdataScr_wb_0),
	.datad(always1),
	.cin(gnd),
	.combout(dataScr_wb),
	.cout());
// synopsys translate_off
defparam \dataScr_wb~0 .lut_mask = 16'hAAF0;
defparam \dataScr_wb~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N28
cycloneive_lcell_comb \dataScr_wb~1 (
// Equation(s):
// dataScr_wb1 = (always1 & (\prif.dataScr_mem [1])) # (!always1 & ((\prif.dataScr_wb [1])))

	.dataa(gnd),
	.datab(prifdataScr_mem_1),
	.datac(prifdataScr_wb_1),
	.datad(always1),
	.cin(gnd),
	.combout(dataScr_wb1),
	.cout());
// synopsys translate_off
defparam \dataScr_wb~1 .lut_mask = 16'hCCF0;
defparam \dataScr_wb~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N2
cycloneive_lcell_comb \pc_wb~0 (
// Equation(s):
// pc_wb = (always1 & ((\prif.pc_mem [1]))) # (!always1 & (\prif.pc_wb [1]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_1),
	.datad(prifpc_mem_1),
	.cin(gnd),
	.combout(pc_wb),
	.cout());
// synopsys translate_off
defparam \pc_wb~0 .lut_mask = 16'hFC30;
defparam \pc_wb~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N20
cycloneive_lcell_comb \rdat2_ex~1 (
// Equation(s):
// rdat2_ex = (ccifiwait_0 & (\prif.rdat2_ex [1])) # (!ccifiwait_0 & ((\rdat2_ex~0_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_1),
	.datad(\rdat2_ex~0_combout ),
	.cin(gnd),
	.combout(rdat2_ex),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~1 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N26
cycloneive_lcell_comb \prif.rs_ex[1]~0 (
// Equation(s):
// prifrs_ex_11 = (\prif.rs_ex[0]~0_combout  & (\prif.rs_ex [1])) # (!\prif.rs_ex[0]~0_combout  & ((\prif.imemload_id [22])))

	.dataa(gnd),
	.datab(prifrs_ex_01),
	.datac(prifrs_ex_1),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(prifrs_ex_11),
	.cout());
// synopsys translate_off
defparam \prif.rs_ex[1]~0 .lut_mask = 16'hF3C0;
defparam \prif.rs_ex[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N16
cycloneive_lcell_comb \prif.rs_ex[0]~1 (
// Equation(s):
// prifrs_ex_02 = (\prif.rs_ex[0]~0_combout  & (\prif.rs_ex [0])) # (!\prif.rs_ex[0]~0_combout  & ((\prif.imemload_id [21])))

	.dataa(gnd),
	.datab(prifrs_ex_01),
	.datac(prifrs_ex_0),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(prifrs_ex_02),
	.cout());
// synopsys translate_off
defparam \prif.rs_ex[0]~1 .lut_mask = 16'hF3C0;
defparam \prif.rs_ex[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N20
cycloneive_lcell_comb \prif.rs_ex[3]~2 (
// Equation(s):
// prifrs_ex_31 = (\prif.rs_ex[0]~0_combout  & (\prif.rs_ex [3])) # (!\prif.rs_ex[0]~0_combout  & ((\prif.imemload_id [24])))

	.dataa(gnd),
	.datab(prifrs_ex_01),
	.datac(prifrs_ex_3),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(prifrs_ex_31),
	.cout());
// synopsys translate_off
defparam \prif.rs_ex[3]~2 .lut_mask = 16'hF3C0;
defparam \prif.rs_ex[3]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N30
cycloneive_lcell_comb \prif.rs_ex[2]~3 (
// Equation(s):
// prifrs_ex_21 = (\prif.rs_ex[0]~0_combout  & (\prif.rs_ex [2])) # (!\prif.rs_ex[0]~0_combout  & ((\prif.imemload_id [23])))

	.dataa(gnd),
	.datab(prifrs_ex_01),
	.datac(prifrs_ex_2),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(prifrs_ex_21),
	.cout());
// synopsys translate_off
defparam \prif.rs_ex[2]~3 .lut_mask = 16'hF3C0;
defparam \prif.rs_ex[2]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y27_N6
cycloneive_lcell_comb \prif.rs_ex[4]~4 (
// Equation(s):
// prifrs_ex_41 = (\prif.rs_ex[0]~0_combout  & (\prif.rs_ex [4])) # (!\prif.rs_ex[0]~0_combout  & ((\prif.imemload_id [25])))

	.dataa(gnd),
	.datab(prifrs_ex_01),
	.datac(prifrs_ex_4),
	.datad(prifimemload_id_25),
	.cin(gnd),
	.combout(prifrs_ex_41),
	.cout());
// synopsys translate_off
defparam \prif.rs_ex[4]~4 .lut_mask = 16'hF3C0;
defparam \prif.rs_ex[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N0
cycloneive_lcell_comb \opcode_mem~0 (
// Equation(s):
// opcode_mem = (exmem_en & (\prif.opcode_ex [1])) # (!exmem_en & ((\prif.opcode_mem [1])))

	.dataa(exmem_en),
	.datab(prifopcode_ex_1),
	.datac(prifopcode_mem_1),
	.datad(gnd),
	.cin(gnd),
	.combout(opcode_mem),
	.cout());
// synopsys translate_off
defparam \opcode_mem~0 .lut_mask = 16'hD8D8;
defparam \opcode_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N6
cycloneive_lcell_comb \opcode_mem~1 (
// Equation(s):
// opcode_mem1 = (exmem_en & (\prif.opcode_ex [0])) # (!exmem_en & ((\prif.opcode_mem [0])))

	.dataa(exmem_en),
	.datab(prifopcode_ex_0),
	.datac(prifopcode_mem_0),
	.datad(gnd),
	.cin(gnd),
	.combout(opcode_mem1),
	.cout());
// synopsys translate_off
defparam \opcode_mem~1 .lut_mask = 16'hD8D8;
defparam \opcode_mem~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N12
cycloneive_lcell_comb \opcode_mem~2 (
// Equation(s):
// opcode_mem2 = (exmem_en & (\prif.opcode_ex [2])) # (!exmem_en & ((\prif.opcode_mem [2])))

	.dataa(prifopcode_ex_2),
	.datab(gnd),
	.datac(prifopcode_mem_2),
	.datad(exmem_en),
	.cin(gnd),
	.combout(opcode_mem2),
	.cout());
// synopsys translate_off
defparam \opcode_mem~2 .lut_mask = 16'hAAF0;
defparam \opcode_mem~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N2
cycloneive_lcell_comb \opcode_mem~3 (
// Equation(s):
// opcode_mem3 = (exmem_en & ((\prif.opcode_ex [3]))) # (!exmem_en & (\prif.opcode_mem [3]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifopcode_mem_3),
	.datad(prifopcode_ex_3),
	.cin(gnd),
	.combout(opcode_mem3),
	.cout());
// synopsys translate_off
defparam \opcode_mem~3 .lut_mask = 16'hFA50;
defparam \opcode_mem~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N24
cycloneive_lcell_comb \opcode_mem~4 (
// Equation(s):
// opcode_mem4 = (exmem_en & ((\prif.opcode_ex [5]))) # (!exmem_en & (\prif.opcode_mem [5]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifopcode_mem_5),
	.datad(prifopcode_ex_5),
	.cin(gnd),
	.combout(opcode_mem4),
	.cout());
// synopsys translate_off
defparam \opcode_mem~4 .lut_mask = 16'hFA50;
defparam \opcode_mem~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N26
cycloneive_lcell_comb \opcode_mem~5 (
// Equation(s):
// opcode_mem5 = (exmem_en & ((\prif.opcode_ex [4]))) # (!exmem_en & (\prif.opcode_mem [4]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifopcode_mem_4),
	.datad(prifopcode_ex_4),
	.cin(gnd),
	.combout(opcode_mem5),
	.cout());
// synopsys translate_off
defparam \opcode_mem~5 .lut_mask = 16'hFA50;
defparam \opcode_mem~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N28
cycloneive_lcell_comb \rdat1_ex~1 (
// Equation(s):
// rdat1_ex = (ccifiwait_0 & (\prif.rdat1_ex [1])) # (!ccifiwait_0 & ((\rdat1_ex~0_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_1),
	.datad(\rdat1_ex~0_combout ),
	.cin(gnd),
	.combout(rdat1_ex),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~1 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N8
cycloneive_lcell_comb \imm_ex~1 (
// Equation(s):
// imm_ex1 = (ccifiwait_0 & (\prif.imm_ex [0])) # (!ccifiwait_0 & ((\prif.imemload_id [0])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifimm_ex_0),
	.datad(prifimemload_id_0),
	.cin(gnd),
	.combout(imm_ex1),
	.cout());
// synopsys translate_off
defparam \imm_ex~1 .lut_mask = 16'hF5A0;
defparam \imm_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N2
cycloneive_lcell_comb \shamt_ex~1 (
// Equation(s):
// shamt_ex1 = (ccifiwait_0 & ((\prif.shamt_ex [0]))) # (!ccifiwait_0 & (\prif.imemload_id [6]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_6),
	.datac(prifshamt_ex_0),
	.datad(gnd),
	.cin(gnd),
	.combout(shamt_ex1),
	.cout());
// synopsys translate_off
defparam \shamt_ex~1 .lut_mask = 16'hE4E4;
defparam \shamt_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N18
cycloneive_lcell_comb \dmemload_wb~1 (
// Equation(s):
// dmemload_wb1 = (always1 & (ramiframload_0)) # (!always1 & ((\prif.dmemload_wb [0])))

	.dataa(ramiframload_0),
	.datab(always1),
	.datac(prifdmemload_wb_0),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemload_wb1),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~1 .lut_mask = 16'hB8B8;
defparam \dmemload_wb~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N20
cycloneive_lcell_comb \dmemaddr_wb~1 (
// Equation(s):
// dmemaddr_wb1 = (always1 & ((prifdmemaddr_0))) # (!always1 & (\prif.dmemaddr_wb [0]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_0),
	.datad(prifdmemaddr_0),
	.cin(gnd),
	.combout(dmemaddr_wb1),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~1 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N0
cycloneive_lcell_comb \pc_wb~1 (
// Equation(s):
// pc_wb1 = (always1 & (\prif.pc_mem [0])) # (!always1 & ((\prif.pc_wb [0])))

	.dataa(prifpc_mem_0),
	.datab(always1),
	.datac(prifpc_wb_0),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_wb1),
	.cout());
// synopsys translate_off
defparam \pc_wb~1 .lut_mask = 16'hB8B8;
defparam \pc_wb~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N16
cycloneive_lcell_comb \rdat2_ex~3 (
// Equation(s):
// rdat2_ex1 = (ccifiwait_0 & (\prif.rdat2_ex [0])) # (!ccifiwait_0 & ((\rdat2_ex~2_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_0),
	.datad(\rdat2_ex~2_combout ),
	.cin(gnd),
	.combout(rdat2_ex1),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~3 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N10
cycloneive_lcell_comb \rdat1_ex~3 (
// Equation(s):
// rdat1_ex1 = (ccifiwait_0 & (\prif.rdat1_ex [0])) # (!ccifiwait_0 & ((\rdat1_ex~2_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_0),
	.datad(\rdat1_ex~2_combout ),
	.cin(gnd),
	.combout(rdat1_ex1),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~3 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N12
cycloneive_lcell_comb \dmemload_wb~2 (
// Equation(s):
// dmemload_wb2 = (always1 & (ramiframload_3)) # (!always1 & ((\prif.dmemload_wb [3])))

	.dataa(ramiframload_3),
	.datab(gnd),
	.datac(prifdmemload_wb_3),
	.datad(always1),
	.cin(gnd),
	.combout(dmemload_wb2),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~2 .lut_mask = 16'hAAF0;
defparam \dmemload_wb~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N26
cycloneive_lcell_comb \dmemaddr_wb~2 (
// Equation(s):
// dmemaddr_wb2 = (always1 & (prifdmemaddr_3)) # (!always1 & ((\prif.dmemaddr_wb [3])))

	.dataa(gnd),
	.datab(prifdmemaddr_3),
	.datac(prifdmemaddr_wb_3),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb2),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~2 .lut_mask = 16'hCCF0;
defparam \dmemaddr_wb~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N10
cycloneive_lcell_comb \pc_wb~2 (
// Equation(s):
// pc_wb2 = (always1 & (\prif.pc_mem [3])) # (!always1 & ((\prif.pc_wb [3])))

	.dataa(prifpc_mem_3),
	.datab(gnd),
	.datac(prifpc_wb_3),
	.datad(always1),
	.cin(gnd),
	.combout(pc_wb2),
	.cout());
// synopsys translate_off
defparam \pc_wb~2 .lut_mask = 16'hAAF0;
defparam \pc_wb~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N0
cycloneive_lcell_comb \rdat2_ex~5 (
// Equation(s):
// rdat2_ex2 = (ccifiwait_0 & (\prif.rdat2_ex [3])) # (!ccifiwait_0 & ((\rdat2_ex~4_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_3),
	.datad(\rdat2_ex~4_combout ),
	.cin(gnd),
	.combout(rdat2_ex2),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~5 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N18
cycloneive_lcell_comb \imm_ex~2 (
// Equation(s):
// imm_ex2 = (ccifiwait_0 & ((\prif.imm_ex [3]))) # (!ccifiwait_0 & (\prif.imemload_id [3]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_3),
	.datac(prifimm_ex_3),
	.datad(gnd),
	.cin(gnd),
	.combout(imm_ex2),
	.cout());
// synopsys translate_off
defparam \imm_ex~2 .lut_mask = 16'hE4E4;
defparam \imm_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N28
cycloneive_lcell_comb \shamt_ex~2 (
// Equation(s):
// shamt_ex2 = (ccifiwait_0 & ((\prif.shamt_ex [3]))) # (!ccifiwait_0 & (\prif.imemload_id [9]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_9),
	.datac(prifshamt_ex_3),
	.datad(gnd),
	.cin(gnd),
	.combout(shamt_ex2),
	.cout());
// synopsys translate_off
defparam \shamt_ex~2 .lut_mask = 16'hE4E4;
defparam \shamt_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N12
cycloneive_lcell_comb \imm_ex~3 (
// Equation(s):
// imm_ex3 = (ccifiwait_0 & (\prif.imm_ex [2])) # (!ccifiwait_0 & ((\prif.imemload_id [2])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifimm_ex_2),
	.datad(prifimemload_id_2),
	.cin(gnd),
	.combout(imm_ex3),
	.cout());
// synopsys translate_off
defparam \imm_ex~3 .lut_mask = 16'hF3C0;
defparam \imm_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N20
cycloneive_lcell_comb \shamt_ex~3 (
// Equation(s):
// shamt_ex3 = (ccifiwait_0 & ((\prif.shamt_ex [2]))) # (!ccifiwait_0 & (\prif.imemload_id [8]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_8),
	.datac(prifshamt_ex_2),
	.datad(gnd),
	.cin(gnd),
	.combout(shamt_ex3),
	.cout());
// synopsys translate_off
defparam \shamt_ex~3 .lut_mask = 16'hE4E4;
defparam \shamt_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N6
cycloneive_lcell_comb \dmemload_wb~3 (
// Equation(s):
// dmemload_wb3 = (always1 & ((ramiframload_2))) # (!always1 & (\prif.dmemload_wb [2]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemload_wb_2),
	.datad(ramiframload_2),
	.cin(gnd),
	.combout(dmemload_wb3),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~3 .lut_mask = 16'hFC30;
defparam \dmemload_wb~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N4
cycloneive_lcell_comb \dmemaddr_wb~3 (
// Equation(s):
// dmemaddr_wb3 = (always1 & ((prifdmemaddr_2))) # (!always1 & (\prif.dmemaddr_wb [2]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_2),
	.datad(prifdmemaddr_2),
	.cin(gnd),
	.combout(dmemaddr_wb3),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~3 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N28
cycloneive_lcell_comb \pc_wb~3 (
// Equation(s):
// pc_wb3 = (always1 & ((\prif.pc_mem [2]))) # (!always1 & (\prif.pc_wb [2]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_2),
	.datad(prifpc_mem_2),
	.cin(gnd),
	.combout(pc_wb3),
	.cout());
// synopsys translate_off
defparam \pc_wb~3 .lut_mask = 16'hFC30;
defparam \pc_wb~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N22
cycloneive_lcell_comb \rdat2_ex~7 (
// Equation(s):
// rdat2_ex3 = (ccifiwait_0 & (\prif.rdat2_ex [2])) # (!ccifiwait_0 & ((\rdat2_ex~6_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_2),
	.datad(\rdat2_ex~6_combout ),
	.cin(gnd),
	.combout(rdat2_ex3),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~7 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N22
cycloneive_lcell_comb \dmemload_wb~4 (
// Equation(s):
// dmemload_wb4 = (always1 & ((ramiframload_4))) # (!always1 & (\prif.dmemload_wb [4]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemload_wb_4),
	.datad(ramiframload_4),
	.cin(gnd),
	.combout(dmemload_wb4),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~4 .lut_mask = 16'hFA50;
defparam \dmemload_wb~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N16
cycloneive_lcell_comb \dmemaddr_wb~4 (
// Equation(s):
// dmemaddr_wb4 = (always1 & (prifdmemaddr_4)) # (!always1 & ((\prif.dmemaddr_wb [4])))

	.dataa(prifdmemaddr_4),
	.datab(gnd),
	.datac(prifdmemaddr_wb_4),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb4),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~4 .lut_mask = 16'hAAF0;
defparam \dmemaddr_wb~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N8
cycloneive_lcell_comb \pc_wb~4 (
// Equation(s):
// pc_wb4 = (always1 & ((\prif.pc_mem [4]))) # (!always1 & (\prif.pc_wb [4]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifpc_wb_4),
	.datad(prifpc_mem_4),
	.cin(gnd),
	.combout(pc_wb4),
	.cout());
// synopsys translate_off
defparam \pc_wb~4 .lut_mask = 16'hFA50;
defparam \pc_wb~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N30
cycloneive_lcell_comb \rdat2_ex~9 (
// Equation(s):
// rdat2_ex4 = (ccifiwait_0 & (\prif.rdat2_ex [4])) # (!ccifiwait_0 & ((\rdat2_ex~8_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_4),
	.datad(\rdat2_ex~8_combout ),
	.cin(gnd),
	.combout(rdat2_ex4),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~9 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N26
cycloneive_lcell_comb \imm_ex~4 (
// Equation(s):
// imm_ex4 = (ccifiwait_0 & (\prif.imm_ex [4])) # (!ccifiwait_0 & ((\prif.imemload_id [4])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifimm_ex_4),
	.datad(prifimemload_id_4),
	.cin(gnd),
	.combout(imm_ex4),
	.cout());
// synopsys translate_off
defparam \imm_ex~4 .lut_mask = 16'hF3C0;
defparam \imm_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N4
cycloneive_lcell_comb \shamt_ex~4 (
// Equation(s):
// shamt_ex4 = (ccifiwait_0 & (\prif.shamt_ex [4])) # (!ccifiwait_0 & ((\prif.imemload_id [10])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifshamt_ex_4),
	.datad(prifimemload_id_10),
	.cin(gnd),
	.combout(shamt_ex4),
	.cout());
// synopsys translate_off
defparam \shamt_ex~4 .lut_mask = 16'hF3C0;
defparam \shamt_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N20
cycloneive_lcell_comb \instr_ex~0 (
// Equation(s):
// instr_ex = (ccifiwait_0 & ((\prif.instr_ex [15]))) # (!ccifiwait_0 & (\prif.imemload_id [15]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_15),
	.datac(prifinstr_ex_15),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_ex),
	.cout());
// synopsys translate_off
defparam \instr_ex~0 .lut_mask = 16'hE4E4;
defparam \instr_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N12
cycloneive_lcell_comb \dmemload_wb~5 (
// Equation(s):
// dmemload_wb5 = (always1 & ((ramiframload_31))) # (!always1 & (\prif.dmemload_wb [31]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemload_wb_31),
	.datad(ramiframload_31),
	.cin(gnd),
	.combout(dmemload_wb5),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~5 .lut_mask = 16'hFA50;
defparam \dmemload_wb~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N26
cycloneive_lcell_comb \imm_wb~0 (
// Equation(s):
// imm_wb = (always1 & (\prif.imm_mem [15])) # (!always1 & ((\prif.imm_wb [15])))

	.dataa(gnd),
	.datab(prifimm_mem_15),
	.datac(prifimm_wb_15),
	.datad(always1),
	.cin(gnd),
	.combout(imm_wb),
	.cout());
// synopsys translate_off
defparam \imm_wb~0 .lut_mask = 16'hCCF0;
defparam \imm_wb~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N16
cycloneive_lcell_comb \dmemaddr_wb~5 (
// Equation(s):
// dmemaddr_wb5 = (always1 & ((prifdmemaddr_31))) # (!always1 & (\prif.dmemaddr_wb [31]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemaddr_wb_31),
	.datad(prifdmemaddr_31),
	.cin(gnd),
	.combout(dmemaddr_wb5),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~5 .lut_mask = 16'hFA50;
defparam \dmemaddr_wb~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N4
cycloneive_lcell_comb \pc_wb~5 (
// Equation(s):
// pc_wb5 = (always1 & ((\prif.pc_mem [31]))) # (!always1 & (\prif.pc_wb [31]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifpc_wb_31),
	.datad(prifpc_mem_31),
	.cin(gnd),
	.combout(pc_wb5),
	.cout());
// synopsys translate_off
defparam \pc_wb~5 .lut_mask = 16'hFA50;
defparam \pc_wb~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y25_N4
cycloneive_lcell_comb \rdat2_ex~11 (
// Equation(s):
// rdat2_ex5 = (ccifiwait_0 & (\prif.rdat2_ex [31])) # (!ccifiwait_0 & ((\rdat2_ex~10_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_31),
	.datad(\rdat2_ex~10_combout ),
	.cin(gnd),
	.combout(rdat2_ex5),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~11 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N22
cycloneive_lcell_comb \imm_mem~0 (
// Equation(s):
// imm_mem = (exmem_en & ((\prif.imm_ex [15]))) # (!exmem_en & (\prif.imm_mem [15]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_15),
	.datad(prifimm_ex_15),
	.cin(gnd),
	.combout(imm_mem),
	.cout());
// synopsys translate_off
defparam \imm_mem~0 .lut_mask = 16'hFA50;
defparam \imm_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N16
cycloneive_lcell_comb \imm_wb~1 (
// Equation(s):
// imm_wb1 = (always1 & (\prif.imm_mem [14])) # (!always1 & ((\prif.imm_wb [14])))

	.dataa(prifimm_mem_14),
	.datab(always1),
	.datac(prifimm_wb_14),
	.datad(gnd),
	.cin(gnd),
	.combout(imm_wb1),
	.cout());
// synopsys translate_off
defparam \imm_wb~1 .lut_mask = 16'hB8B8;
defparam \imm_wb~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N30
cycloneive_lcell_comb \dmemload_wb~6 (
// Equation(s):
// dmemload_wb6 = (always1 & (ramiframload_30)) # (!always1 & ((\prif.dmemload_wb [30])))

	.dataa(always1),
	.datab(ramiframload_30),
	.datac(prifdmemload_wb_30),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemload_wb6),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~6 .lut_mask = 16'hD8D8;
defparam \dmemload_wb~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N20
cycloneive_lcell_comb \dmemaddr_wb~6 (
// Equation(s):
// dmemaddr_wb6 = (always1 & ((prifdmemaddr_30))) # (!always1 & (\prif.dmemaddr_wb [30]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_30),
	.datad(prifdmemaddr_30),
	.cin(gnd),
	.combout(dmemaddr_wb6),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~6 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N4
cycloneive_lcell_comb \pc_wb~6 (
// Equation(s):
// pc_wb6 = (always1 & ((\prif.pc_mem [30]))) # (!always1 & (\prif.pc_wb [30]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_30),
	.datad(prifpc_mem_30),
	.cin(gnd),
	.combout(pc_wb6),
	.cout());
// synopsys translate_off
defparam \pc_wb~6 .lut_mask = 16'hFC30;
defparam \pc_wb~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N0
cycloneive_lcell_comb \rdat2_ex~13 (
// Equation(s):
// rdat2_ex6 = (ccifiwait_0 & (\prif.rdat2_ex [30])) # (!ccifiwait_0 & ((\rdat2_ex~12_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_30),
	.datad(\rdat2_ex~12_combout ),
	.cin(gnd),
	.combout(rdat2_ex6),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~13 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N26
cycloneive_lcell_comb \imm_mem~1 (
// Equation(s):
// imm_mem1 = (exmem_en & ((\prif.imm_ex [14]))) # (!exmem_en & (\prif.imm_mem [14]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_14),
	.datad(prifimm_ex_14),
	.cin(gnd),
	.combout(imm_mem1),
	.cout());
// synopsys translate_off
defparam \imm_mem~1 .lut_mask = 16'hFA50;
defparam \imm_mem~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N22
cycloneive_lcell_comb \dmemload_wb~7 (
// Equation(s):
// dmemload_wb7 = (always1 & ((ramiframload_29))) # (!always1 & (\prif.dmemload_wb [29]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemload_wb_29),
	.datad(ramiframload_29),
	.cin(gnd),
	.combout(dmemload_wb7),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~7 .lut_mask = 16'hFC30;
defparam \dmemload_wb~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N12
cycloneive_lcell_comb \imm_wb~2 (
// Equation(s):
// imm_wb2 = (always1 & ((\prif.imm_mem [13]))) # (!always1 & (\prif.imm_wb [13]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifimm_wb_13),
	.datad(prifimm_mem_13),
	.cin(gnd),
	.combout(imm_wb2),
	.cout());
// synopsys translate_off
defparam \imm_wb~2 .lut_mask = 16'hFC30;
defparam \imm_wb~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N10
cycloneive_lcell_comb \dmemaddr_wb~7 (
// Equation(s):
// dmemaddr_wb7 = (always1 & ((prifdmemaddr_29))) # (!always1 & (\prif.dmemaddr_wb [29]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_29),
	.datad(prifdmemaddr_29),
	.cin(gnd),
	.combout(dmemaddr_wb7),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~7 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N14
cycloneive_lcell_comb \pc_wb~7 (
// Equation(s):
// pc_wb7 = (always1 & ((\prif.pc_mem [29]))) # (!always1 & (\prif.pc_wb [29]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_29),
	.datad(prifpc_mem_29),
	.cin(gnd),
	.combout(pc_wb7),
	.cout());
// synopsys translate_off
defparam \pc_wb~7 .lut_mask = 16'hFC30;
defparam \pc_wb~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N6
cycloneive_lcell_comb \rdat2_ex~15 (
// Equation(s):
// rdat2_ex7 = (ccifiwait_0 & (\prif.rdat2_ex [29])) # (!ccifiwait_0 & ((\rdat2_ex~14_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_29),
	.datad(\rdat2_ex~14_combout ),
	.cin(gnd),
	.combout(rdat2_ex7),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~15 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N2
cycloneive_lcell_comb \imm_mem~2 (
// Equation(s):
// imm_mem2 = (exmem_en & ((\prif.imm_ex [13]))) # (!exmem_en & (\prif.imm_mem [13]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_13),
	.datad(prifimm_ex_13),
	.cin(gnd),
	.combout(imm_mem2),
	.cout());
// synopsys translate_off
defparam \imm_mem~2 .lut_mask = 16'hFA50;
defparam \imm_mem~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N16
cycloneive_lcell_comb \imm_ex~5 (
// Equation(s):
// imm_ex5 = (ccifiwait_0 & (\prif.imm_ex [5])) # (!ccifiwait_0 & ((\prif.imemload_id [5])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifimm_ex_5),
	.datad(prifimemload_id_5),
	.cin(gnd),
	.combout(imm_ex5),
	.cout());
// synopsys translate_off
defparam \imm_ex~5 .lut_mask = 16'hF3C0;
defparam \imm_ex~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N20
cycloneive_lcell_comb \dmemload_wb~8 (
// Equation(s):
// dmemload_wb8 = (always1 & ((ramiframload_5))) # (!always1 & (\prif.dmemload_wb [5]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemload_wb_5),
	.datad(ramiframload_5),
	.cin(gnd),
	.combout(dmemload_wb8),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~8 .lut_mask = 16'hFA50;
defparam \dmemload_wb~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N22
cycloneive_lcell_comb \dmemaddr_wb~8 (
// Equation(s):
// dmemaddr_wb8 = (always1 & ((prifdmemaddr_5))) # (!always1 & (\prif.dmemaddr_wb [5]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemaddr_wb_5),
	.datad(prifdmemaddr_5),
	.cin(gnd),
	.combout(dmemaddr_wb8),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~8 .lut_mask = 16'hFA50;
defparam \dmemaddr_wb~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N12
cycloneive_lcell_comb \pc_wb~8 (
// Equation(s):
// pc_wb8 = (always1 & ((\prif.pc_mem [5]))) # (!always1 & (\prif.pc_wb [5]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifpc_wb_5),
	.datad(prifpc_mem_5),
	.cin(gnd),
	.combout(pc_wb8),
	.cout());
// synopsys translate_off
defparam \pc_wb~8 .lut_mask = 16'hFA50;
defparam \pc_wb~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N4
cycloneive_lcell_comb \rdat2_ex~17 (
// Equation(s):
// rdat2_ex8 = (ccifiwait_0 & ((\prif.rdat2_ex [5]))) # (!ccifiwait_0 & (\rdat2_ex~16_combout ))

	.dataa(\rdat2_ex~16_combout ),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_5),
	.datad(gnd),
	.cin(gnd),
	.combout(rdat2_ex8),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~17 .lut_mask = 16'hE2E2;
defparam \rdat2_ex~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N22
cycloneive_lcell_comb \imm_ex~6 (
// Equation(s):
// imm_ex6 = (ccifiwait_0 & ((\prif.imm_ex [15]))) # (!ccifiwait_0 & (\prif.imemload_id [15]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_15),
	.datac(prifimm_ex_15),
	.datad(gnd),
	.cin(gnd),
	.combout(imm_ex6),
	.cout());
// synopsys translate_off
defparam \imm_ex~6 .lut_mask = 16'hE4E4;
defparam \imm_ex~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N30
cycloneive_lcell_comb \dmemload_wb~9 (
// Equation(s):
// dmemload_wb9 = (always1 & ((ramiframload_15))) # (!always1 & (\prif.dmemload_wb [15]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemload_wb_15),
	.datad(ramiframload_15),
	.cin(gnd),
	.combout(dmemload_wb9),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~9 .lut_mask = 16'hFA50;
defparam \dmemload_wb~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N2
cycloneive_lcell_comb \dmemaddr_wb~9 (
// Equation(s):
// dmemaddr_wb9 = (always1 & (prifdmemaddr_15)) # (!always1 & ((\prif.dmemaddr_wb [15])))

	.dataa(always1),
	.datab(prifdmemaddr_15),
	.datac(prifdmemaddr_wb_15),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemaddr_wb9),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~9 .lut_mask = 16'hD8D8;
defparam \dmemaddr_wb~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N26
cycloneive_lcell_comb \pc_wb~9 (
// Equation(s):
// pc_wb9 = (always1 & (\prif.pc_mem [15])) # (!always1 & ((\prif.pc_wb [15])))

	.dataa(prifpc_mem_15),
	.datab(gnd),
	.datac(prifpc_wb_15),
	.datad(always1),
	.cin(gnd),
	.combout(pc_wb9),
	.cout());
// synopsys translate_off
defparam \pc_wb~9 .lut_mask = 16'hAAF0;
defparam \pc_wb~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N28
cycloneive_lcell_comb \rdat2_ex~19 (
// Equation(s):
// rdat2_ex9 = (ccifiwait_0 & (\prif.rdat2_ex [15])) # (!ccifiwait_0 & ((\rdat2_ex~18_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_15),
	.datad(\rdat2_ex~18_combout ),
	.cin(gnd),
	.combout(rdat2_ex9),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~19 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N16
cycloneive_lcell_comb \imm_ex~7 (
// Equation(s):
// imm_ex7 = (ccifiwait_0 & (\prif.imm_ex [14])) # (!ccifiwait_0 & ((\prif.imemload_id [14])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifimm_ex_14),
	.datad(prifimemload_id_14),
	.cin(gnd),
	.combout(imm_ex7),
	.cout());
// synopsys translate_off
defparam \imm_ex~7 .lut_mask = 16'hF5A0;
defparam \imm_ex~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N22
cycloneive_lcell_comb \dmemload_wb~10 (
// Equation(s):
// dmemload_wb10 = (always1 & (ramiframload_14)) # (!always1 & ((\prif.dmemload_wb [14])))

	.dataa(ramiframload_14),
	.datab(gnd),
	.datac(prifdmemload_wb_14),
	.datad(always1),
	.cin(gnd),
	.combout(dmemload_wb10),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~10 .lut_mask = 16'hAAF0;
defparam \dmemload_wb~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N24
cycloneive_lcell_comb \dmemaddr_wb~10 (
// Equation(s):
// dmemaddr_wb10 = (always1 & (prifdmemaddr_14)) # (!always1 & ((\prif.dmemaddr_wb [14])))

	.dataa(gnd),
	.datab(prifdmemaddr_14),
	.datac(prifdmemaddr_wb_14),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb10),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~10 .lut_mask = 16'hCCF0;
defparam \dmemaddr_wb~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N28
cycloneive_lcell_comb \pc_wb~10 (
// Equation(s):
// pc_wb10 = (always1 & ((\prif.pc_mem [14]))) # (!always1 & (\prif.pc_wb [14]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_14),
	.datad(prifpc_mem_14),
	.cin(gnd),
	.combout(pc_wb10),
	.cout());
// synopsys translate_off
defparam \pc_wb~10 .lut_mask = 16'hFC30;
defparam \pc_wb~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N20
cycloneive_lcell_comb \rdat2_ex~21 (
// Equation(s):
// rdat2_ex10 = (ccifiwait_0 & (\prif.rdat2_ex [14])) # (!ccifiwait_0 & ((\rdat2_ex~20_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_14),
	.datad(\rdat2_ex~20_combout ),
	.cin(gnd),
	.combout(rdat2_ex10),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~21 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N28
cycloneive_lcell_comb \imm_ex~8 (
// Equation(s):
// imm_ex8 = (ccifiwait_0 & (\prif.imm_ex [13])) # (!ccifiwait_0 & ((\prif.imemload_id [13])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifimm_ex_13),
	.datad(prifimemload_id_13),
	.cin(gnd),
	.combout(imm_ex8),
	.cout());
// synopsys translate_off
defparam \imm_ex~8 .lut_mask = 16'hF5A0;
defparam \imm_ex~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N12
cycloneive_lcell_comb \dmemload_wb~11 (
// Equation(s):
// dmemload_wb11 = (always1 & (ramiframload_13)) # (!always1 & ((\prif.dmemload_wb [13])))

	.dataa(ramiframload_13),
	.datab(gnd),
	.datac(prifdmemload_wb_13),
	.datad(always1),
	.cin(gnd),
	.combout(dmemload_wb11),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~11 .lut_mask = 16'hAAF0;
defparam \dmemload_wb~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N2
cycloneive_lcell_comb \dmemaddr_wb~11 (
// Equation(s):
// dmemaddr_wb11 = (always1 & (prifdmemaddr_13)) # (!always1 & ((\prif.dmemaddr_wb [13])))

	.dataa(prifdmemaddr_13),
	.datab(gnd),
	.datac(prifdmemaddr_wb_13),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb11),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~11 .lut_mask = 16'hAAF0;
defparam \dmemaddr_wb~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N22
cycloneive_lcell_comb \pc_wb~11 (
// Equation(s):
// pc_wb11 = (always1 & ((\prif.pc_mem [13]))) # (!always1 & (\prif.pc_wb [13]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_13),
	.datad(prifpc_mem_13),
	.cin(gnd),
	.combout(pc_wb11),
	.cout());
// synopsys translate_off
defparam \pc_wb~11 .lut_mask = 16'hFC30;
defparam \pc_wb~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N26
cycloneive_lcell_comb \rdat2_ex~23 (
// Equation(s):
// rdat2_ex11 = (ccifiwait_0 & (\prif.rdat2_ex [13])) # (!ccifiwait_0 & ((\rdat2_ex~22_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_13),
	.datad(\rdat2_ex~22_combout ),
	.cin(gnd),
	.combout(rdat2_ex11),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~23 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N0
cycloneive_lcell_comb \imm_ex~9 (
// Equation(s):
// imm_ex9 = (ccifiwait_0 & (\prif.imm_ex [12])) # (!ccifiwait_0 & ((\prif.imemload_id [12])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifimm_ex_12),
	.datad(prifimemload_id_12),
	.cin(gnd),
	.combout(imm_ex9),
	.cout());
// synopsys translate_off
defparam \imm_ex~9 .lut_mask = 16'hF3C0;
defparam \imm_ex~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N20
cycloneive_lcell_comb \dmemload_wb~12 (
// Equation(s):
// dmemload_wb12 = (always1 & (ramiframload_12)) # (!always1 & ((\prif.dmemload_wb [12])))

	.dataa(always1),
	.datab(ramiframload_12),
	.datac(prifdmemload_wb_12),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemload_wb12),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~12 .lut_mask = 16'hD8D8;
defparam \dmemload_wb~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N30
cycloneive_lcell_comb \dmemaddr_wb~12 (
// Equation(s):
// dmemaddr_wb12 = (always1 & (prifdmemaddr_12)) # (!always1 & ((\prif.dmemaddr_wb [12])))

	.dataa(always1),
	.datab(prifdmemaddr_12),
	.datac(prifdmemaddr_wb_12),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemaddr_wb12),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~12 .lut_mask = 16'hD8D8;
defparam \dmemaddr_wb~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N26
cycloneive_lcell_comb \pc_wb~12 (
// Equation(s):
// pc_wb12 = (always1 & (\prif.pc_mem [12])) # (!always1 & ((\prif.pc_wb [12])))

	.dataa(always1),
	.datab(prifpc_mem_12),
	.datac(prifpc_wb_12),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_wb12),
	.cout());
// synopsys translate_off
defparam \pc_wb~12 .lut_mask = 16'hD8D8;
defparam \pc_wb~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N10
cycloneive_lcell_comb \rdat2_ex~25 (
// Equation(s):
// rdat2_ex12 = (ccifiwait_0 & (\prif.rdat2_ex [12])) # (!ccifiwait_0 & ((\rdat2_ex~24_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_12),
	.datad(\rdat2_ex~24_combout ),
	.cin(gnd),
	.combout(rdat2_ex12),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~25 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N22
cycloneive_lcell_comb \imm_ex~10 (
// Equation(s):
// imm_ex10 = (ccifiwait_0 & ((\prif.imm_ex [11]))) # (!ccifiwait_0 & (\prif.imemload_id [11]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_11),
	.datac(prifimm_ex_11),
	.datad(gnd),
	.cin(gnd),
	.combout(imm_ex10),
	.cout());
// synopsys translate_off
defparam \imm_ex~10 .lut_mask = 16'hE4E4;
defparam \imm_ex~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N6
cycloneive_lcell_comb \dmemload_wb~13 (
// Equation(s):
// dmemload_wb13 = (always1 & (ramiframload_11)) # (!always1 & ((\prif.dmemload_wb [11])))

	.dataa(ramiframload_11),
	.datab(always1),
	.datac(prifdmemload_wb_11),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemload_wb13),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~13 .lut_mask = 16'hB8B8;
defparam \dmemload_wb~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N28
cycloneive_lcell_comb \dmemaddr_wb~13 (
// Equation(s):
// dmemaddr_wb13 = (always1 & ((prifdmemaddr_11))) # (!always1 & (\prif.dmemaddr_wb [11]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_11),
	.datad(prifdmemaddr_11),
	.cin(gnd),
	.combout(dmemaddr_wb13),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~13 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N8
cycloneive_lcell_comb \pc_wb~13 (
// Equation(s):
// pc_wb13 = (always1 & ((\prif.pc_mem [11]))) # (!always1 & (\prif.pc_wb [11]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_11),
	.datad(prifpc_mem_11),
	.cin(gnd),
	.combout(pc_wb13),
	.cout());
// synopsys translate_off
defparam \pc_wb~13 .lut_mask = 16'hFC30;
defparam \pc_wb~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N26
cycloneive_lcell_comb \rdat2_ex~27 (
// Equation(s):
// rdat2_ex13 = (ccifiwait_0 & (\prif.rdat2_ex [11])) # (!ccifiwait_0 & ((\rdat2_ex~26_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_11),
	.datad(\rdat2_ex~26_combout ),
	.cin(gnd),
	.combout(rdat2_ex13),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~27 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N10
cycloneive_lcell_comb \imm_ex~11 (
// Equation(s):
// imm_ex11 = (ccifiwait_0 & (\prif.imm_ex [10])) # (!ccifiwait_0 & ((\prif.imemload_id [10])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifimm_ex_10),
	.datad(prifimemload_id_10),
	.cin(gnd),
	.combout(imm_ex11),
	.cout());
// synopsys translate_off
defparam \imm_ex~11 .lut_mask = 16'hF3C0;
defparam \imm_ex~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N8
cycloneive_lcell_comb \dmemload_wb~14 (
// Equation(s):
// dmemload_wb14 = (always1 & (ramiframload_10)) # (!always1 & ((\prif.dmemload_wb [10])))

	.dataa(ramiframload_10),
	.datab(always1),
	.datac(prifdmemload_wb_10),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemload_wb14),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~14 .lut_mask = 16'hB8B8;
defparam \dmemload_wb~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N30
cycloneive_lcell_comb \dmemaddr_wb~14 (
// Equation(s):
// dmemaddr_wb14 = (always1 & ((prifdmemaddr_10))) # (!always1 & (\prif.dmemaddr_wb [10]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_10),
	.datad(prifdmemaddr_10),
	.cin(gnd),
	.combout(dmemaddr_wb14),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~14 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N22
cycloneive_lcell_comb \pc_wb~14 (
// Equation(s):
// pc_wb14 = (always1 & ((\prif.pc_mem [10]))) # (!always1 & (\prif.pc_wb [10]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_10),
	.datad(prifpc_mem_10),
	.cin(gnd),
	.combout(pc_wb14),
	.cout());
// synopsys translate_off
defparam \pc_wb~14 .lut_mask = 16'hFC30;
defparam \pc_wb~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N0
cycloneive_lcell_comb \rdat2_ex~29 (
// Equation(s):
// rdat2_ex14 = (ccifiwait_0 & (\prif.rdat2_ex [10])) # (!ccifiwait_0 & ((\rdat2_ex~28_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_10),
	.datad(\rdat2_ex~28_combout ),
	.cin(gnd),
	.combout(rdat2_ex14),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~29 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N10
cycloneive_lcell_comb \imm_ex~12 (
// Equation(s):
// imm_ex12 = (ccifiwait_0 & (\prif.imm_ex [9])) # (!ccifiwait_0 & ((\prif.imemload_id [9])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifimm_ex_9),
	.datad(prifimemload_id_9),
	.cin(gnd),
	.combout(imm_ex12),
	.cout());
// synopsys translate_off
defparam \imm_ex~12 .lut_mask = 16'hF3C0;
defparam \imm_ex~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N28
cycloneive_lcell_comb \dmemload_wb~15 (
// Equation(s):
// dmemload_wb15 = (always1 & (ramiframload_9)) # (!always1 & ((\prif.dmemload_wb [9])))

	.dataa(always1),
	.datab(ramiframload_9),
	.datac(prifdmemload_wb_9),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemload_wb15),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~15 .lut_mask = 16'hD8D8;
defparam \dmemload_wb~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N6
cycloneive_lcell_comb \dmemaddr_wb~15 (
// Equation(s):
// dmemaddr_wb15 = (always1 & ((prifdmemaddr_9))) # (!always1 & (\prif.dmemaddr_wb [9]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_9),
	.datad(prifdmemaddr_9),
	.cin(gnd),
	.combout(dmemaddr_wb15),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~15 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N22
cycloneive_lcell_comb \pc_wb~15 (
// Equation(s):
// pc_wb15 = (always1 & ((\prif.pc_mem [9]))) # (!always1 & (\prif.pc_wb [9]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifpc_wb_9),
	.datad(prifpc_mem_9),
	.cin(gnd),
	.combout(pc_wb15),
	.cout());
// synopsys translate_off
defparam \pc_wb~15 .lut_mask = 16'hFA50;
defparam \pc_wb~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N4
cycloneive_lcell_comb \rdat2_ex~31 (
// Equation(s):
// rdat2_ex15 = (ccifiwait_0 & (\prif.rdat2_ex [9])) # (!ccifiwait_0 & ((\rdat2_ex~30_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_9),
	.datad(\rdat2_ex~30_combout ),
	.cin(gnd),
	.combout(rdat2_ex15),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~31 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N4
cycloneive_lcell_comb \imm_ex~13 (
// Equation(s):
// imm_ex13 = (ccifiwait_0 & (\prif.imm_ex [6])) # (!ccifiwait_0 & ((\prif.imemload_id [6])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifimm_ex_6),
	.datad(prifimemload_id_6),
	.cin(gnd),
	.combout(imm_ex13),
	.cout());
// synopsys translate_off
defparam \imm_ex~13 .lut_mask = 16'hF5A0;
defparam \imm_ex~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N2
cycloneive_lcell_comb \dmemload_wb~16 (
// Equation(s):
// dmemload_wb16 = (always1 & (ramiframload_6)) # (!always1 & ((\prif.dmemload_wb [6])))

	.dataa(ramiframload_6),
	.datab(always1),
	.datac(prifdmemload_wb_6),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemload_wb16),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~16 .lut_mask = 16'hB8B8;
defparam \dmemload_wb~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N4
cycloneive_lcell_comb \dmemaddr_wb~16 (
// Equation(s):
// dmemaddr_wb16 = (always1 & ((prifdmemaddr_6))) # (!always1 & (\prif.dmemaddr_wb [6]))

	.dataa(prifdmemaddr_wb_6),
	.datab(prifdmemaddr_6),
	.datac(always1),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemaddr_wb16),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~16 .lut_mask = 16'hCACA;
defparam \dmemaddr_wb~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N24
cycloneive_lcell_comb \pc_wb~16 (
// Equation(s):
// pc_wb16 = (always1 & ((\prif.pc_mem [6]))) # (!always1 & (\prif.pc_wb [6]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifpc_wb_6),
	.datad(prifpc_mem_6),
	.cin(gnd),
	.combout(pc_wb16),
	.cout());
// synopsys translate_off
defparam \pc_wb~16 .lut_mask = 16'hFA50;
defparam \pc_wb~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N30
cycloneive_lcell_comb \rdat2_ex~33 (
// Equation(s):
// rdat2_ex16 = (ccifiwait_0 & (\prif.rdat2_ex [6])) # (!ccifiwait_0 & ((\rdat2_ex~32_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_6),
	.datad(\rdat2_ex~32_combout ),
	.cin(gnd),
	.combout(rdat2_ex16),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~33 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N16
cycloneive_lcell_comb \dmemload_wb~17 (
// Equation(s):
// dmemload_wb17 = (always1 & ((ramiframload_27))) # (!always1 & (\prif.dmemload_wb [27]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemload_wb_27),
	.datad(ramiframload_27),
	.cin(gnd),
	.combout(dmemload_wb17),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~17 .lut_mask = 16'hFA50;
defparam \dmemload_wb~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N10
cycloneive_lcell_comb \imm_wb~3 (
// Equation(s):
// imm_wb3 = (always1 & (\prif.imm_mem [11])) # (!always1 & ((\prif.imm_wb [11])))

	.dataa(prifimm_mem_11),
	.datab(gnd),
	.datac(prifimm_wb_11),
	.datad(always1),
	.cin(gnd),
	.combout(imm_wb3),
	.cout());
// synopsys translate_off
defparam \imm_wb~3 .lut_mask = 16'hAAF0;
defparam \imm_wb~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N0
cycloneive_lcell_comb \dmemaddr_wb~17 (
// Equation(s):
// dmemaddr_wb17 = (always1 & ((prifdmemaddr_27))) # (!always1 & (\prif.dmemaddr_wb [27]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemaddr_wb_27),
	.datad(prifdmemaddr_27),
	.cin(gnd),
	.combout(dmemaddr_wb17),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~17 .lut_mask = 16'hFA50;
defparam \dmemaddr_wb~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N12
cycloneive_lcell_comb \pc_wb~17 (
// Equation(s):
// pc_wb17 = (always1 & ((\prif.pc_mem [27]))) # (!always1 & (\prif.pc_wb [27]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifpc_wb_27),
	.datad(prifpc_mem_27),
	.cin(gnd),
	.combout(pc_wb17),
	.cout());
// synopsys translate_off
defparam \pc_wb~17 .lut_mask = 16'hFA50;
defparam \pc_wb~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N20
cycloneive_lcell_comb \rdat2_ex~35 (
// Equation(s):
// rdat2_ex17 = (ccifiwait_0 & (\prif.rdat2_ex [27])) # (!ccifiwait_0 & ((\rdat2_ex~34_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_27),
	.datad(\rdat2_ex~34_combout ),
	.cin(gnd),
	.combout(rdat2_ex17),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~35 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N30
cycloneive_lcell_comb \imm_mem~3 (
// Equation(s):
// imm_mem3 = (exmem_en & (\prif.imm_ex [11])) # (!exmem_en & ((\prif.imm_mem [11])))

	.dataa(exmem_en),
	.datab(prifimm_ex_11),
	.datac(prifimm_mem_11),
	.datad(gnd),
	.cin(gnd),
	.combout(imm_mem3),
	.cout());
// synopsys translate_off
defparam \imm_mem~3 .lut_mask = 16'hD8D8;
defparam \imm_mem~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N4
cycloneive_lcell_comb \dmemload_wb~18 (
// Equation(s):
// dmemload_wb18 = (always1 & ((ramiframload_23))) # (!always1 & (\prif.dmemload_wb [23]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemload_wb_23),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(dmemload_wb18),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~18 .lut_mask = 16'hFC30;
defparam \dmemload_wb~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N14
cycloneive_lcell_comb \imm_wb~4 (
// Equation(s):
// imm_wb4 = (always1 & ((\prif.imm_mem [7]))) # (!always1 & (\prif.imm_wb [7]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifimm_wb_7),
	.datad(prifimm_mem_7),
	.cin(gnd),
	.combout(imm_wb4),
	.cout());
// synopsys translate_off
defparam \imm_wb~4 .lut_mask = 16'hFC30;
defparam \imm_wb~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N24
cycloneive_lcell_comb \dmemaddr_wb~18 (
// Equation(s):
// dmemaddr_wb18 = (always1 & (prifdmemaddr_23)) # (!always1 & ((\prif.dmemaddr_wb [23])))

	.dataa(prifdmemaddr_23),
	.datab(gnd),
	.datac(prifdmemaddr_wb_23),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb18),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~18 .lut_mask = 16'hAAF0;
defparam \dmemaddr_wb~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N12
cycloneive_lcell_comb \pc_wb~18 (
// Equation(s):
// pc_wb18 = (always1 & ((\prif.pc_mem [23]))) # (!always1 & (\prif.pc_wb [23]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_23),
	.datad(prifpc_mem_23),
	.cin(gnd),
	.combout(pc_wb18),
	.cout());
// synopsys translate_off
defparam \pc_wb~18 .lut_mask = 16'hFC30;
defparam \pc_wb~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N26
cycloneive_lcell_comb \rdat2_ex~37 (
// Equation(s):
// rdat2_ex18 = (ccifiwait_0 & (\prif.rdat2_ex [23])) # (!ccifiwait_0 & ((\rdat2_ex~36_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_23),
	.datad(\rdat2_ex~36_combout ),
	.cin(gnd),
	.combout(rdat2_ex18),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~37 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N16
cycloneive_lcell_comb \imm_mem~4 (
// Equation(s):
// imm_mem4 = (exmem_en & ((\prif.imm_ex [7]))) # (!exmem_en & (\prif.imm_mem [7]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifimm_mem_7),
	.datad(prifimm_ex_7),
	.cin(gnd),
	.combout(imm_mem4),
	.cout());
// synopsys translate_off
defparam \imm_mem~4 .lut_mask = 16'hFC30;
defparam \imm_mem~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N18
cycloneive_lcell_comb \imm_wb~5 (
// Equation(s):
// imm_wb5 = (always1 & (\prif.imm_mem [2])) # (!always1 & ((\prif.imm_wb [2])))

	.dataa(gnd),
	.datab(prifimm_mem_2),
	.datac(prifimm_wb_2),
	.datad(always1),
	.cin(gnd),
	.combout(imm_wb5),
	.cout());
// synopsys translate_off
defparam \imm_wb~5 .lut_mask = 16'hCCF0;
defparam \imm_wb~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N0
cycloneive_lcell_comb \dmemload_wb~19 (
// Equation(s):
// dmemload_wb19 = (always1 & (ramiframload_18)) # (!always1 & ((\prif.dmemload_wb [18])))

	.dataa(gnd),
	.datab(ramiframload_18),
	.datac(prifdmemload_wb_18),
	.datad(always1),
	.cin(gnd),
	.combout(dmemload_wb19),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~19 .lut_mask = 16'hCCF0;
defparam \dmemload_wb~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N2
cycloneive_lcell_comb \dmemaddr_wb~19 (
// Equation(s):
// dmemaddr_wb19 = (always1 & (prifdmemaddr_18)) # (!always1 & ((\prif.dmemaddr_wb [18])))

	.dataa(prifdmemaddr_18),
	.datab(gnd),
	.datac(prifdmemaddr_wb_18),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb19),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~19 .lut_mask = 16'hAAF0;
defparam \dmemaddr_wb~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N30
cycloneive_lcell_comb \pc_wb~19 (
// Equation(s):
// pc_wb19 = (always1 & (\prif.pc_mem [18])) # (!always1 & ((\prif.pc_wb [18])))

	.dataa(prifpc_mem_18),
	.datab(gnd),
	.datac(prifpc_wb_18),
	.datad(always1),
	.cin(gnd),
	.combout(pc_wb19),
	.cout());
// synopsys translate_off
defparam \pc_wb~19 .lut_mask = 16'hAAF0;
defparam \pc_wb~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N8
cycloneive_lcell_comb \rdat2_ex~39 (
// Equation(s):
// rdat2_ex19 = (ccifiwait_0 & (\prif.rdat2_ex [18])) # (!ccifiwait_0 & ((\rdat2_ex~38_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_18),
	.datad(\rdat2_ex~38_combout ),
	.cin(gnd),
	.combout(rdat2_ex19),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~39 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N8
cycloneive_lcell_comb \imm_mem~5 (
// Equation(s):
// imm_mem5 = (exmem_en & ((\prif.imm_ex [2]))) # (!exmem_en & (\prif.imm_mem [2]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifimm_mem_2),
	.datad(prifimm_ex_2),
	.cin(gnd),
	.combout(imm_mem5),
	.cout());
// synopsys translate_off
defparam \imm_mem~5 .lut_mask = 16'hFC30;
defparam \imm_mem~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N26
cycloneive_lcell_comb \imm_wb~6 (
// Equation(s):
// imm_wb6 = (always1 & ((\prif.imm_mem [8]))) # (!always1 & (\prif.imm_wb [8]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifimm_wb_8),
	.datad(prifimm_mem_8),
	.cin(gnd),
	.combout(imm_wb6),
	.cout());
// synopsys translate_off
defparam \imm_wb~6 .lut_mask = 16'hFA50;
defparam \imm_wb~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N16
cycloneive_lcell_comb \dmemload_wb~20 (
// Equation(s):
// dmemload_wb20 = (always1 & ((ramiframload_24))) # (!always1 & (\prif.dmemload_wb [24]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemload_wb_24),
	.datad(ramiframload_24),
	.cin(gnd),
	.combout(dmemload_wb20),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~20 .lut_mask = 16'hFA50;
defparam \dmemload_wb~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N22
cycloneive_lcell_comb \dmemaddr_wb~20 (
// Equation(s):
// dmemaddr_wb20 = (always1 & ((prifdmemaddr_24))) # (!always1 & (\prif.dmemaddr_wb [24]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemaddr_wb_24),
	.datad(prifdmemaddr_24),
	.cin(gnd),
	.combout(dmemaddr_wb20),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~20 .lut_mask = 16'hFA50;
defparam \dmemaddr_wb~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N18
cycloneive_lcell_comb \pc_wb~20 (
// Equation(s):
// pc_wb20 = (always1 & ((\prif.pc_mem [24]))) # (!always1 & (\prif.pc_wb [24]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifpc_wb_24),
	.datad(prifpc_mem_24),
	.cin(gnd),
	.combout(pc_wb20),
	.cout());
// synopsys translate_off
defparam \pc_wb~20 .lut_mask = 16'hFA50;
defparam \pc_wb~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N18
cycloneive_lcell_comb \rdat2_ex~41 (
// Equation(s):
// rdat2_ex20 = (ccifiwait_0 & (\prif.rdat2_ex [24])) # (!ccifiwait_0 & ((\rdat2_ex~40_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_24),
	.datad(\rdat2_ex~40_combout ),
	.cin(gnd),
	.combout(rdat2_ex20),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~41 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N12
cycloneive_lcell_comb \imm_mem~6 (
// Equation(s):
// imm_mem6 = (exmem_en & (\prif.imm_ex [8])) # (!exmem_en & ((\prif.imm_mem [8])))

	.dataa(prifimm_ex_8),
	.datab(gnd),
	.datac(prifimm_mem_8),
	.datad(exmem_en),
	.cin(gnd),
	.combout(imm_mem6),
	.cout());
// synopsys translate_off
defparam \imm_mem~6 .lut_mask = 16'hAAF0;
defparam \imm_mem~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N0
cycloneive_lcell_comb \imm_wb~7 (
// Equation(s):
// imm_wb7 = (always1 & ((\prif.imm_mem [0]))) # (!always1 & (\prif.imm_wb [0]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifimm_wb_0),
	.datad(prifimm_mem_0),
	.cin(gnd),
	.combout(imm_wb7),
	.cout());
// synopsys translate_off
defparam \imm_wb~7 .lut_mask = 16'hFC30;
defparam \imm_wb~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N4
cycloneive_lcell_comb \dmemload_wb~21 (
// Equation(s):
// dmemload_wb21 = (always1 & ((ramiframload_16))) # (!always1 & (\prif.dmemload_wb [16]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemload_wb_16),
	.datad(ramiframload_16),
	.cin(gnd),
	.combout(dmemload_wb21),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~21 .lut_mask = 16'hFA50;
defparam \dmemload_wb~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N26
cycloneive_lcell_comb \dmemaddr_wb~21 (
// Equation(s):
// dmemaddr_wb21 = (always1 & ((prifdmemaddr_16))) # (!always1 & (\prif.dmemaddr_wb [16]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemaddr_wb_16),
	.datad(prifdmemaddr_16),
	.cin(gnd),
	.combout(dmemaddr_wb21),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~21 .lut_mask = 16'hFA50;
defparam \dmemaddr_wb~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N2
cycloneive_lcell_comb \pc_wb~21 (
// Equation(s):
// pc_wb21 = (always1 & ((\prif.pc_mem [16]))) # (!always1 & (\prif.pc_wb [16]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_16),
	.datad(prifpc_mem_16),
	.cin(gnd),
	.combout(pc_wb21),
	.cout());
// synopsys translate_off
defparam \pc_wb~21 .lut_mask = 16'hFC30;
defparam \pc_wb~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N4
cycloneive_lcell_comb \rdat2_ex~43 (
// Equation(s):
// rdat2_ex21 = (ccifiwait_0 & (\prif.rdat2_ex [16])) # (!ccifiwait_0 & ((\rdat2_ex~42_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_16),
	.datad(\rdat2_ex~42_combout ),
	.cin(gnd),
	.combout(rdat2_ex21),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~43 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N2
cycloneive_lcell_comb \imm_mem~7 (
// Equation(s):
// imm_mem7 = (exmem_en & ((\prif.imm_ex [0]))) # (!exmem_en & (\prif.imm_mem [0]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_0),
	.datad(prifimm_ex_0),
	.cin(gnd),
	.combout(imm_mem7),
	.cout());
// synopsys translate_off
defparam \imm_mem~7 .lut_mask = 16'hFA50;
defparam \imm_mem~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N8
cycloneive_lcell_comb \dmemload_wb~22 (
// Equation(s):
// dmemload_wb22 = (always1 & ((ramiframload_19))) # (!always1 & (\prif.dmemload_wb [19]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemload_wb_19),
	.datad(ramiframload_19),
	.cin(gnd),
	.combout(dmemload_wb22),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~22 .lut_mask = 16'hFC30;
defparam \dmemload_wb~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N22
cycloneive_lcell_comb \imm_wb~8 (
// Equation(s):
// imm_wb8 = (always1 & (\prif.imm_mem [3])) # (!always1 & ((\prif.imm_wb [3])))

	.dataa(prifimm_mem_3),
	.datab(always1),
	.datac(prifimm_wb_3),
	.datad(gnd),
	.cin(gnd),
	.combout(imm_wb8),
	.cout());
// synopsys translate_off
defparam \imm_wb~8 .lut_mask = 16'hB8B8;
defparam \imm_wb~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N20
cycloneive_lcell_comb \dmemaddr_wb~22 (
// Equation(s):
// dmemaddr_wb22 = (always1 & ((prifdmemaddr_19))) # (!always1 & (\prif.dmemaddr_wb [19]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_19),
	.datad(prifdmemaddr_19),
	.cin(gnd),
	.combout(dmemaddr_wb22),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~22 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N16
cycloneive_lcell_comb \pc_wb~22 (
// Equation(s):
// pc_wb22 = (always1 & ((\prif.pc_mem [19]))) # (!always1 & (\prif.pc_wb [19]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_19),
	.datad(prifpc_mem_19),
	.cin(gnd),
	.combout(pc_wb22),
	.cout());
// synopsys translate_off
defparam \pc_wb~22 .lut_mask = 16'hFC30;
defparam \pc_wb~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N26
cycloneive_lcell_comb \rdat2_ex~45 (
// Equation(s):
// rdat2_ex22 = (ccifiwait_0 & (\prif.rdat2_ex [19])) # (!ccifiwait_0 & ((\rdat2_ex~44_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_19),
	.datad(\rdat2_ex~44_combout ),
	.cin(gnd),
	.combout(rdat2_ex22),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~45 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y29_N26
cycloneive_lcell_comb \imm_mem~8 (
// Equation(s):
// imm_mem8 = (exmem_en & ((\prif.imm_ex [3]))) # (!exmem_en & (\prif.imm_mem [3]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_3),
	.datad(prifimm_ex_3),
	.cin(gnd),
	.combout(imm_mem8),
	.cout());
// synopsys translate_off
defparam \imm_mem~8 .lut_mask = 16'hFA50;
defparam \imm_mem~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N18
cycloneive_lcell_comb \dmemload_wb~23 (
// Equation(s):
// dmemload_wb23 = (always1 & ((ramiframload_17))) # (!always1 & (\prif.dmemload_wb [17]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifdmemload_wb_17),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(dmemload_wb23),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~23 .lut_mask = 16'hFA50;
defparam \dmemload_wb~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N0
cycloneive_lcell_comb \imm_wb~9 (
// Equation(s):
// imm_wb9 = (always1 & ((\prif.imm_mem [1]))) # (!always1 & (\prif.imm_wb [1]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifimm_wb_1),
	.datad(prifimm_mem_1),
	.cin(gnd),
	.combout(imm_wb9),
	.cout());
// synopsys translate_off
defparam \imm_wb~9 .lut_mask = 16'hFA50;
defparam \imm_wb~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N22
cycloneive_lcell_comb \dmemaddr_wb~23 (
// Equation(s):
// dmemaddr_wb23 = (always1 & (prifdmemaddr_17)) # (!always1 & ((\prif.dmemaddr_wb [17])))

	.dataa(prifdmemaddr_17),
	.datab(gnd),
	.datac(prifdmemaddr_wb_17),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb23),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~23 .lut_mask = 16'hAAF0;
defparam \dmemaddr_wb~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N22
cycloneive_lcell_comb \pc_wb~23 (
// Equation(s):
// pc_wb23 = (always1 & ((\prif.pc_mem [17]))) # (!always1 & (\prif.pc_wb [17]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifpc_wb_17),
	.datad(prifpc_mem_17),
	.cin(gnd),
	.combout(pc_wb23),
	.cout());
// synopsys translate_off
defparam \pc_wb~23 .lut_mask = 16'hFA50;
defparam \pc_wb~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N8
cycloneive_lcell_comb \rdat2_ex~47 (
// Equation(s):
// rdat2_ex23 = (ccifiwait_0 & (\prif.rdat2_ex [17])) # (!ccifiwait_0 & ((\rdat2_ex~46_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_17),
	.datad(\rdat2_ex~46_combout ),
	.cin(gnd),
	.combout(rdat2_ex23),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~47 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N28
cycloneive_lcell_comb \imm_mem~9 (
// Equation(s):
// imm_mem9 = (exmem_en & ((\prif.imm_ex [1]))) # (!exmem_en & (\prif.imm_mem [1]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_1),
	.datad(prifimm_ex_1),
	.cin(gnd),
	.combout(imm_mem9),
	.cout());
// synopsys translate_off
defparam \imm_mem~9 .lut_mask = 16'hFA50;
defparam \imm_mem~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N20
cycloneive_lcell_comb \dmemload_wb~24 (
// Equation(s):
// dmemload_wb24 = (always1 & (ramiframload_21)) # (!always1 & ((\prif.dmemload_wb [21])))

	.dataa(gnd),
	.datab(ramiframload_21),
	.datac(prifdmemload_wb_21),
	.datad(always1),
	.cin(gnd),
	.combout(dmemload_wb24),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~24 .lut_mask = 16'hCCF0;
defparam \dmemload_wb~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N0
cycloneive_lcell_comb \imm_wb~10 (
// Equation(s):
// imm_wb10 = (always1 & ((\prif.imm_mem [5]))) # (!always1 & (\prif.imm_wb [5]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifimm_wb_5),
	.datad(prifimm_mem_5),
	.cin(gnd),
	.combout(imm_wb10),
	.cout());
// synopsys translate_off
defparam \imm_wb~10 .lut_mask = 16'hFC30;
defparam \imm_wb~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N26
cycloneive_lcell_comb \dmemaddr_wb~24 (
// Equation(s):
// dmemaddr_wb24 = (always1 & ((prifdmemaddr_21))) # (!always1 & (\prif.dmemaddr_wb [21]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_21),
	.datad(prifdmemaddr_21),
	.cin(gnd),
	.combout(dmemaddr_wb24),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~24 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N18
cycloneive_lcell_comb \pc_wb~24 (
// Equation(s):
// pc_wb24 = (always1 & ((\prif.pc_mem [21]))) # (!always1 & (\prif.pc_wb [21]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_21),
	.datad(prifpc_mem_21),
	.cin(gnd),
	.combout(pc_wb24),
	.cout());
// synopsys translate_off
defparam \pc_wb~24 .lut_mask = 16'hFC30;
defparam \pc_wb~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N20
cycloneive_lcell_comb \rdat2_ex~49 (
// Equation(s):
// rdat2_ex24 = (ccifiwait_0 & (\prif.rdat2_ex [21])) # (!ccifiwait_0 & ((\rdat2_ex~48_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_21),
	.datad(\rdat2_ex~48_combout ),
	.cin(gnd),
	.combout(rdat2_ex24),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~49 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N4
cycloneive_lcell_comb \imm_mem~10 (
// Equation(s):
// imm_mem10 = (exmem_en & ((\prif.imm_ex [5]))) # (!exmem_en & (\prif.imm_mem [5]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_5),
	.datad(prifimm_ex_5),
	.cin(gnd),
	.combout(imm_mem10),
	.cout());
// synopsys translate_off
defparam \imm_mem~10 .lut_mask = 16'hFA50;
defparam \imm_mem~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N26
cycloneive_lcell_comb \imm_wb~11 (
// Equation(s):
// imm_wb11 = (always1 & ((\prif.imm_mem [4]))) # (!always1 & (\prif.imm_wb [4]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifimm_wb_4),
	.datad(prifimm_mem_4),
	.cin(gnd),
	.combout(imm_wb11),
	.cout());
// synopsys translate_off
defparam \imm_wb~11 .lut_mask = 16'hFA50;
defparam \imm_wb~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N12
cycloneive_lcell_comb \dmemload_wb~25 (
// Equation(s):
// dmemload_wb25 = (always1 & (ramiframload_20)) # (!always1 & ((\prif.dmemload_wb [20])))

	.dataa(always1),
	.datab(ramiframload_20),
	.datac(prifdmemload_wb_20),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemload_wb25),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~25 .lut_mask = 16'hD8D8;
defparam \dmemload_wb~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N18
cycloneive_lcell_comb \dmemaddr_wb~25 (
// Equation(s):
// dmemaddr_wb25 = (always1 & (prifdmemaddr_20)) # (!always1 & ((\prif.dmemaddr_wb [20])))

	.dataa(always1),
	.datab(prifdmemaddr_20),
	.datac(prifdmemaddr_wb_20),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemaddr_wb25),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~25 .lut_mask = 16'hD8D8;
defparam \dmemaddr_wb~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N30
cycloneive_lcell_comb \pc_wb~25 (
// Equation(s):
// pc_wb25 = (always1 & (\prif.pc_mem [20])) # (!always1 & ((\prif.pc_wb [20])))

	.dataa(always1),
	.datab(prifpc_mem_20),
	.datac(prifpc_wb_20),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_wb25),
	.cout());
// synopsys translate_off
defparam \pc_wb~25 .lut_mask = 16'hD8D8;
defparam \pc_wb~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N4
cycloneive_lcell_comb \rdat2_ex~51 (
// Equation(s):
// rdat2_ex25 = (ccifiwait_0 & (\prif.rdat2_ex [20])) # (!ccifiwait_0 & ((\rdat2_ex~50_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_20),
	.datad(\rdat2_ex~50_combout ),
	.cin(gnd),
	.combout(rdat2_ex25),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~51 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N30
cycloneive_lcell_comb \imm_mem~11 (
// Equation(s):
// imm_mem11 = (exmem_en & ((\prif.imm_ex [4]))) # (!exmem_en & (\prif.imm_mem [4]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_4),
	.datad(prifimm_ex_4),
	.cin(gnd),
	.combout(imm_mem11),
	.cout());
// synopsys translate_off
defparam \imm_mem~11 .lut_mask = 16'hFA50;
defparam \imm_mem~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N0
cycloneive_lcell_comb \imm_wb~12 (
// Equation(s):
// imm_wb12 = (always1 & ((\prif.imm_mem [12]))) # (!always1 & (\prif.imm_wb [12]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifimm_wb_12),
	.datad(prifimm_mem_12),
	.cin(gnd),
	.combout(imm_wb12),
	.cout());
// synopsys translate_off
defparam \imm_wb~12 .lut_mask = 16'hFC30;
defparam \imm_wb~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N22
cycloneive_lcell_comb \dmemload_wb~26 (
// Equation(s):
// dmemload_wb26 = (always1 & ((ramiframload_28))) # (!always1 & (\prif.dmemload_wb [28]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemload_wb_28),
	.datad(ramiframload_28),
	.cin(gnd),
	.combout(dmemload_wb26),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~26 .lut_mask = 16'hFC30;
defparam \dmemload_wb~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N4
cycloneive_lcell_comb \dmemaddr_wb~26 (
// Equation(s):
// dmemaddr_wb26 = (always1 & (prifdmemaddr_28)) # (!always1 & ((\prif.dmemaddr_wb [28])))

	.dataa(gnd),
	.datab(prifdmemaddr_28),
	.datac(prifdmemaddr_wb_28),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb26),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~26 .lut_mask = 16'hCCF0;
defparam \dmemaddr_wb~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N12
cycloneive_lcell_comb \pc_wb~26 (
// Equation(s):
// pc_wb26 = (always1 & (\prif.pc_mem [28])) # (!always1 & ((\prif.pc_wb [28])))

	.dataa(prifpc_mem_28),
	.datab(gnd),
	.datac(prifpc_wb_28),
	.datad(always1),
	.cin(gnd),
	.combout(pc_wb26),
	.cout());
// synopsys translate_off
defparam \pc_wb~26 .lut_mask = 16'hAAF0;
defparam \pc_wb~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N24
cycloneive_lcell_comb \rdat2_ex~53 (
// Equation(s):
// rdat2_ex26 = (ccifiwait_0 & (\prif.rdat2_ex [28])) # (!ccifiwait_0 & ((\rdat2_ex~52_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat2_ex_28),
	.datad(\rdat2_ex~52_combout ),
	.cin(gnd),
	.combout(rdat2_ex26),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~53 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N8
cycloneive_lcell_comb \imm_mem~12 (
// Equation(s):
// imm_mem12 = (exmem_en & ((\prif.imm_ex [12]))) # (!exmem_en & (\prif.imm_mem [12]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_12),
	.datad(prifimm_ex_12),
	.cin(gnd),
	.combout(imm_mem12),
	.cout());
// synopsys translate_off
defparam \imm_mem~12 .lut_mask = 16'hFA50;
defparam \imm_mem~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N14
cycloneive_lcell_comb \imm_wb~13 (
// Equation(s):
// imm_wb13 = (always1 & (\prif.imm_mem [10])) # (!always1 & ((\prif.imm_wb [10])))

	.dataa(prifimm_mem_10),
	.datab(always1),
	.datac(prifimm_wb_10),
	.datad(gnd),
	.cin(gnd),
	.combout(imm_wb13),
	.cout());
// synopsys translate_off
defparam \imm_wb~13 .lut_mask = 16'hB8B8;
defparam \imm_wb~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N28
cycloneive_lcell_comb \dmemload_wb~27 (
// Equation(s):
// dmemload_wb27 = (always1 & ((ramiframload_26))) # (!always1 & (\prif.dmemload_wb [26]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemload_wb_26),
	.datad(ramiframload_26),
	.cin(gnd),
	.combout(dmemload_wb27),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~27 .lut_mask = 16'hFC30;
defparam \dmemload_wb~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N10
cycloneive_lcell_comb \dmemaddr_wb~27 (
// Equation(s):
// dmemaddr_wb27 = (always1 & ((prifdmemaddr_26))) # (!always1 & (\prif.dmemaddr_wb [26]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifdmemaddr_wb_26),
	.datad(prifdmemaddr_26),
	.cin(gnd),
	.combout(dmemaddr_wb27),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~27 .lut_mask = 16'hFC30;
defparam \dmemaddr_wb~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N6
cycloneive_lcell_comb \pc_wb~27 (
// Equation(s):
// pc_wb27 = (always1 & ((\prif.pc_mem [26]))) # (!always1 & (\prif.pc_wb [26]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_26),
	.datad(prifpc_mem_26),
	.cin(gnd),
	.combout(pc_wb27),
	.cout());
// synopsys translate_off
defparam \pc_wb~27 .lut_mask = 16'hFC30;
defparam \pc_wb~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N8
cycloneive_lcell_comb \rdat2_ex~55 (
// Equation(s):
// rdat2_ex27 = (ccifiwait_0 & (\prif.rdat2_ex [26])) # (!ccifiwait_0 & ((\rdat2_ex~54_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_26),
	.datad(\rdat2_ex~54_combout ),
	.cin(gnd),
	.combout(rdat2_ex27),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~55 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N26
cycloneive_lcell_comb \imm_mem~13 (
// Equation(s):
// imm_mem13 = (exmem_en & (\prif.imm_ex [10])) # (!exmem_en & ((\prif.imm_mem [10])))

	.dataa(prifimm_ex_10),
	.datab(exmem_en),
	.datac(prifimm_mem_10),
	.datad(gnd),
	.cin(gnd),
	.combout(imm_mem13),
	.cout());
// synopsys translate_off
defparam \imm_mem~13 .lut_mask = 16'hB8B8;
defparam \imm_mem~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N14
cycloneive_lcell_comb \imm_ex~14 (
// Equation(s):
// imm_ex14 = (ccifiwait_0 & (\prif.imm_ex [8])) # (!ccifiwait_0 & ((\prif.imemload_id [8])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifimm_ex_8),
	.datad(prifimemload_id_8),
	.cin(gnd),
	.combout(imm_ex14),
	.cout());
// synopsys translate_off
defparam \imm_ex~14 .lut_mask = 16'hF5A0;
defparam \imm_ex~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N30
cycloneive_lcell_comb \dmemload_wb~28 (
// Equation(s):
// dmemload_wb28 = (always1 & (ramiframload_8)) # (!always1 & ((\prif.dmemload_wb [8])))

	.dataa(gnd),
	.datab(ramiframload_8),
	.datac(prifdmemload_wb_8),
	.datad(always1),
	.cin(gnd),
	.combout(dmemload_wb28),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~28 .lut_mask = 16'hCCF0;
defparam \dmemload_wb~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N2
cycloneive_lcell_comb \dmemaddr_wb~28 (
// Equation(s):
// dmemaddr_wb28 = (always1 & (prifdmemaddr_8)) # (!always1 & ((\prif.dmemaddr_wb [8])))

	.dataa(gnd),
	.datab(prifdmemaddr_8),
	.datac(prifdmemaddr_wb_8),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb28),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~28 .lut_mask = 16'hCCF0;
defparam \dmemaddr_wb~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N16
cycloneive_lcell_comb \pc_wb~28 (
// Equation(s):
// pc_wb28 = (always1 & ((\prif.pc_mem [8]))) # (!always1 & (\prif.pc_wb [8]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_8),
	.datad(prifpc_mem_8),
	.cin(gnd),
	.combout(pc_wb28),
	.cout());
// synopsys translate_off
defparam \pc_wb~28 .lut_mask = 16'hFC30;
defparam \pc_wb~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N30
cycloneive_lcell_comb \rdat2_ex~57 (
// Equation(s):
// rdat2_ex28 = (ccifiwait_0 & (\prif.rdat2_ex [8])) # (!ccifiwait_0 & ((\rdat2_ex~56_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_8),
	.datad(\rdat2_ex~56_combout ),
	.cin(gnd),
	.combout(rdat2_ex28),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~57 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N10
cycloneive_lcell_comb \imm_ex~15 (
// Equation(s):
// imm_ex15 = (ccifiwait_0 & ((\prif.imm_ex [7]))) # (!ccifiwait_0 & (\prif.imemload_id [7]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_7),
	.datac(prifimm_ex_7),
	.datad(gnd),
	.cin(gnd),
	.combout(imm_ex15),
	.cout());
// synopsys translate_off
defparam \imm_ex~15 .lut_mask = 16'hE4E4;
defparam \imm_ex~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N8
cycloneive_lcell_comb \dmemload_wb~29 (
// Equation(s):
// dmemload_wb29 = (always1 & (ramiframload_7)) # (!always1 & ((\prif.dmemload_wb [7])))

	.dataa(gnd),
	.datab(ramiframload_7),
	.datac(prifdmemload_wb_7),
	.datad(always1),
	.cin(gnd),
	.combout(dmemload_wb29),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~29 .lut_mask = 16'hCCF0;
defparam \dmemload_wb~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y29_N10
cycloneive_lcell_comb \dmemaddr_wb~29 (
// Equation(s):
// dmemaddr_wb29 = (always1 & (prifdmemaddr_7)) # (!always1 & ((\prif.dmemaddr_wb [7])))

	.dataa(gnd),
	.datab(prifdmemaddr_7),
	.datac(prifdmemaddr_wb_7),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb29),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~29 .lut_mask = 16'hCCF0;
defparam \dmemaddr_wb~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N18
cycloneive_lcell_comb \pc_wb~29 (
// Equation(s):
// pc_wb29 = (always1 & ((\prif.pc_mem [7]))) # (!always1 & (\prif.pc_wb [7]))

	.dataa(always1),
	.datab(gnd),
	.datac(prifpc_wb_7),
	.datad(prifpc_mem_7),
	.cin(gnd),
	.combout(pc_wb29),
	.cout());
// synopsys translate_off
defparam \pc_wb~29 .lut_mask = 16'hFA50;
defparam \pc_wb~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N16
cycloneive_lcell_comb \rdat2_ex~59 (
// Equation(s):
// rdat2_ex29 = (ccifiwait_0 & (\prif.rdat2_ex [7])) # (!ccifiwait_0 & ((\rdat2_ex~58_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_7),
	.datad(\rdat2_ex~58_combout ),
	.cin(gnd),
	.combout(rdat2_ex29),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~59 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N8
cycloneive_lcell_comb \imm_wb~14 (
// Equation(s):
// imm_wb14 = (always1 & ((\prif.imm_mem [6]))) # (!always1 & (\prif.imm_wb [6]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifimm_wb_6),
	.datad(prifimm_mem_6),
	.cin(gnd),
	.combout(imm_wb14),
	.cout());
// synopsys translate_off
defparam \imm_wb~14 .lut_mask = 16'hFC30;
defparam \imm_wb~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N30
cycloneive_lcell_comb \dmemload_wb~30 (
// Equation(s):
// dmemload_wb30 = (always1 & (ramiframload_22)) # (!always1 & ((\prif.dmemload_wb [22])))

	.dataa(ramiframload_22),
	.datab(gnd),
	.datac(prifdmemload_wb_22),
	.datad(always1),
	.cin(gnd),
	.combout(dmemload_wb30),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~30 .lut_mask = 16'hAAF0;
defparam \dmemload_wb~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N28
cycloneive_lcell_comb \dmemaddr_wb~30 (
// Equation(s):
// dmemaddr_wb30 = (always1 & (prifdmemaddr_22)) # (!always1 & ((\prif.dmemaddr_wb [22])))

	.dataa(gnd),
	.datab(prifdmemaddr_22),
	.datac(prifdmemaddr_wb_22),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb30),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~30 .lut_mask = 16'hCCF0;
defparam \dmemaddr_wb~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y27_N20
cycloneive_lcell_comb \pc_wb~30 (
// Equation(s):
// pc_wb30 = (always1 & ((\prif.pc_mem [22]))) # (!always1 & (\prif.pc_wb [22]))

	.dataa(gnd),
	.datab(always1),
	.datac(prifpc_wb_22),
	.datad(prifpc_mem_22),
	.cin(gnd),
	.combout(pc_wb30),
	.cout());
// synopsys translate_off
defparam \pc_wb~30 .lut_mask = 16'hFC30;
defparam \pc_wb~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N12
cycloneive_lcell_comb \rdat2_ex~61 (
// Equation(s):
// rdat2_ex30 = (ccifiwait_0 & (\prif.rdat2_ex [22])) # (!ccifiwait_0 & ((\rdat2_ex~60_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_22),
	.datad(\rdat2_ex~60_combout ),
	.cin(gnd),
	.combout(rdat2_ex30),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~61 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y26_N0
cycloneive_lcell_comb \imm_mem~14 (
// Equation(s):
// imm_mem14 = (exmem_en & ((\prif.imm_ex [6]))) # (!exmem_en & (\prif.imm_mem [6]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifimm_mem_6),
	.datad(prifimm_ex_6),
	.cin(gnd),
	.combout(imm_mem14),
	.cout());
// synopsys translate_off
defparam \imm_mem~14 .lut_mask = 16'hFA50;
defparam \imm_mem~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N12
cycloneive_lcell_comb \dmemload_wb~31 (
// Equation(s):
// dmemload_wb31 = (always1 & (ramiframload_25)) # (!always1 & ((\prif.dmemload_wb [25])))

	.dataa(gnd),
	.datab(ramiframload_25),
	.datac(prifdmemload_wb_25),
	.datad(always1),
	.cin(gnd),
	.combout(dmemload_wb31),
	.cout());
// synopsys translate_off
defparam \dmemload_wb~31 .lut_mask = 16'hCCF0;
defparam \dmemload_wb~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N26
cycloneive_lcell_comb \imm_wb~15 (
// Equation(s):
// imm_wb15 = (always1 & (\prif.imm_mem [9])) # (!always1 & ((\prif.imm_wb [9])))

	.dataa(gnd),
	.datab(prifimm_mem_9),
	.datac(prifimm_wb_9),
	.datad(always1),
	.cin(gnd),
	.combout(imm_wb15),
	.cout());
// synopsys translate_off
defparam \imm_wb~15 .lut_mask = 16'hCCF0;
defparam \imm_wb~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N16
cycloneive_lcell_comb \dmemaddr_wb~31 (
// Equation(s):
// dmemaddr_wb31 = (always1 & (prifdmemaddr_25)) # (!always1 & ((\prif.dmemaddr_wb [25])))

	.dataa(gnd),
	.datab(prifdmemaddr_25),
	.datac(prifdmemaddr_wb_25),
	.datad(always1),
	.cin(gnd),
	.combout(dmemaddr_wb31),
	.cout());
// synopsys translate_off
defparam \dmemaddr_wb~31 .lut_mask = 16'hCCF0;
defparam \dmemaddr_wb~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N8
cycloneive_lcell_comb \pc_wb~31 (
// Equation(s):
// pc_wb31 = (always1 & (\prif.pc_mem [25])) # (!always1 & ((\prif.pc_wb [25])))

	.dataa(gnd),
	.datab(prifpc_mem_25),
	.datac(prifpc_wb_25),
	.datad(always1),
	.cin(gnd),
	.combout(pc_wb31),
	.cout());
// synopsys translate_off
defparam \pc_wb~31 .lut_mask = 16'hCCF0;
defparam \pc_wb~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N24
cycloneive_lcell_comb \rdat2_ex~63 (
// Equation(s):
// rdat2_ex31 = (ccifiwait_0 & (\prif.rdat2_ex [25])) # (!ccifiwait_0 & ((\rdat2_ex~62_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat2_ex_25),
	.datad(\rdat2_ex~62_combout ),
	.cin(gnd),
	.combout(rdat2_ex31),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~63 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y28_N24
cycloneive_lcell_comb \imm_mem~15 (
// Equation(s):
// imm_mem15 = (exmem_en & (\prif.imm_ex [9])) # (!exmem_en & ((\prif.imm_mem [9])))

	.dataa(gnd),
	.datab(prifimm_ex_9),
	.datac(prifimm_mem_9),
	.datad(exmem_en),
	.cin(gnd),
	.combout(imm_mem15),
	.cout());
// synopsys translate_off
defparam \imm_mem~15 .lut_mask = 16'hCCF0;
defparam \imm_mem~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N18
cycloneive_lcell_comb \ALUOP_ex~2 (
// Equation(s):
// ALUOP_ex1 = (!flush_idex & ((ccifiwait_0 & (\prif.ALUOP_ex [2])) # (!ccifiwait_0 & ((!\ALUOP_ex~1_combout )))))

	.dataa(flush_idex),
	.datab(ccifiwait_0),
	.datac(prifALUOP_ex_2),
	.datad(\ALUOP_ex~1_combout ),
	.cin(gnd),
	.combout(ALUOP_ex1),
	.cout());
// synopsys translate_off
defparam \ALUOP_ex~2 .lut_mask = 16'h4051;
defparam \ALUOP_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y25_N30
cycloneive_lcell_comb \ALUOP_ex~3 (
// Equation(s):
// ALUOP_ex2 = (!flush_idex & ((ccifiwait_0 & ((\prif.ALUOP_ex [1]))) # (!ccifiwait_0 & (!Selector21))))

	.dataa(Selector21),
	.datab(flush_idex),
	.datac(prifALUOP_ex_1),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(ALUOP_ex2),
	.cout());
// synopsys translate_off
defparam \ALUOP_ex~3 .lut_mask = 16'h3011;
defparam \ALUOP_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N8
cycloneive_lcell_comb \rdat1_ex~5 (
// Equation(s):
// rdat1_ex2 = (ccifiwait_0 & (\prif.rdat1_ex [2])) # (!ccifiwait_0 & ((\rdat1_ex~4_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_2),
	.datad(\rdat1_ex~4_combout ),
	.cin(gnd),
	.combout(rdat1_ex2),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~5 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N0
cycloneive_lcell_comb \rdat1_ex~7 (
// Equation(s):
// rdat1_ex3 = (ccifiwait_0 & (\prif.rdat1_ex [4])) # (!ccifiwait_0 & ((\rdat1_ex~6_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_4),
	.datad(\rdat1_ex~6_combout ),
	.cin(gnd),
	.combout(rdat1_ex3),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~7 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N30
cycloneive_lcell_comb \rdat1_ex~9 (
// Equation(s):
// rdat1_ex4 = (ccifiwait_0 & (\prif.rdat1_ex [3])) # (!ccifiwait_0 & ((\rdat1_ex~8_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_3),
	.datad(\rdat1_ex~8_combout ),
	.cin(gnd),
	.combout(rdat1_ex4),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~9 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N30
cycloneive_lcell_comb \rdat1_ex~11 (
// Equation(s):
// rdat1_ex5 = (ccifiwait_0 & (\prif.rdat1_ex [8])) # (!ccifiwait_0 & ((\rdat1_ex~10_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_8),
	.datad(\rdat1_ex~10_combout ),
	.cin(gnd),
	.combout(rdat1_ex5),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~11 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N30
cycloneive_lcell_comb \rdat1_ex~13 (
// Equation(s):
// rdat1_ex6 = (ccifiwait_0 & (\prif.rdat1_ex [7])) # (!ccifiwait_0 & ((\rdat1_ex~12_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_7),
	.datad(\rdat1_ex~12_combout ),
	.cin(gnd),
	.combout(rdat1_ex6),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~13 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N0
cycloneive_lcell_comb \rdat1_ex~15 (
// Equation(s):
// rdat1_ex7 = (ccifiwait_0 & (\prif.rdat1_ex [6])) # (!ccifiwait_0 & ((\rdat1_ex~14_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_6),
	.datad(\rdat1_ex~14_combout ),
	.cin(gnd),
	.combout(rdat1_ex7),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~15 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N4
cycloneive_lcell_comb \rdat1_ex~17 (
// Equation(s):
// rdat1_ex8 = (ccifiwait_0 & (\prif.rdat1_ex [5])) # (!ccifiwait_0 & ((\rdat1_ex~16_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_5),
	.datad(\rdat1_ex~16_combout ),
	.cin(gnd),
	.combout(rdat1_ex8),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~17 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N22
cycloneive_lcell_comb \rdat1_ex~19 (
// Equation(s):
// rdat1_ex9 = (ccifiwait_0 & (\prif.rdat1_ex [16])) # (!ccifiwait_0 & ((\rdat1_ex~18_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_16),
	.datad(\rdat1_ex~18_combout ),
	.cin(gnd),
	.combout(rdat1_ex9),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~19 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N14
cycloneive_lcell_comb \rdat1_ex~21 (
// Equation(s):
// rdat1_ex10 = (ccifiwait_0 & (\prif.rdat1_ex [15])) # (!ccifiwait_0 & ((\rdat1_ex~20_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_15),
	.datad(\rdat1_ex~20_combout ),
	.cin(gnd),
	.combout(rdat1_ex10),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~21 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N28
cycloneive_lcell_comb \rdat1_ex~23 (
// Equation(s):
// rdat1_ex11 = (ccifiwait_0 & (\prif.rdat1_ex [14])) # (!ccifiwait_0 & ((\rdat1_ex~22_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_14),
	.datad(\rdat1_ex~22_combout ),
	.cin(gnd),
	.combout(rdat1_ex11),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~23 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y26_N20
cycloneive_lcell_comb \rdat1_ex~25 (
// Equation(s):
// rdat1_ex12 = (ccifiwait_0 & (\prif.rdat1_ex [13])) # (!ccifiwait_0 & ((\rdat1_ex~24_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_13),
	.datad(\rdat1_ex~24_combout ),
	.cin(gnd),
	.combout(rdat1_ex12),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~25 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N22
cycloneive_lcell_comb \rdat1_ex~27 (
// Equation(s):
// rdat1_ex13 = (ccifiwait_0 & (\prif.rdat1_ex [11])) # (!ccifiwait_0 & ((\rdat1_ex~26_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_11),
	.datad(\rdat1_ex~26_combout ),
	.cin(gnd),
	.combout(rdat1_ex13),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~27 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N12
cycloneive_lcell_comb \rdat1_ex~29 (
// Equation(s):
// rdat1_ex14 = (ccifiwait_0 & (\prif.rdat1_ex [12])) # (!ccifiwait_0 & ((\rdat1_ex~28_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_12),
	.datad(\rdat1_ex~28_combout ),
	.cin(gnd),
	.combout(rdat1_ex14),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~29 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N22
cycloneive_lcell_comb \rdat1_ex~31 (
// Equation(s):
// rdat1_ex15 = (ccifiwait_0 & (\prif.rdat1_ex [10])) # (!ccifiwait_0 & ((\rdat1_ex~30_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_10),
	.datad(\rdat1_ex~30_combout ),
	.cin(gnd),
	.combout(rdat1_ex15),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~31 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y26_N26
cycloneive_lcell_comb \rdat1_ex~33 (
// Equation(s):
// rdat1_ex16 = (ccifiwait_0 & (\prif.rdat1_ex [9])) # (!ccifiwait_0 & ((\rdat1_ex~32_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_9),
	.datad(\rdat1_ex~32_combout ),
	.cin(gnd),
	.combout(rdat1_ex16),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~33 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N28
cycloneive_lcell_comb \rdat1_ex~35 (
// Equation(s):
// rdat1_ex17 = (ccifiwait_0 & (\prif.rdat1_ex [18])) # (!ccifiwait_0 & ((\rdat1_ex~34_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_18),
	.datad(\rdat1_ex~34_combout ),
	.cin(gnd),
	.combout(rdat1_ex17),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~35 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N14
cycloneive_lcell_comb \rdat1_ex~37 (
// Equation(s):
// rdat1_ex18 = (ccifiwait_0 & (\prif.rdat1_ex [17])) # (!ccifiwait_0 & ((\rdat1_ex~36_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_17),
	.datad(\rdat1_ex~36_combout ),
	.cin(gnd),
	.combout(rdat1_ex18),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~37 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N6
cycloneive_lcell_comb \rdat1_ex~39 (
// Equation(s):
// rdat1_ex19 = (ccifiwait_0 & (\prif.rdat1_ex [20])) # (!ccifiwait_0 & ((\rdat1_ex~38_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_20),
	.datad(\rdat1_ex~38_combout ),
	.cin(gnd),
	.combout(rdat1_ex19),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~39 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N8
cycloneive_lcell_comb \rdat1_ex~41 (
// Equation(s):
// rdat1_ex20 = (ccifiwait_0 & (\prif.rdat1_ex [19])) # (!ccifiwait_0 & ((\rdat1_ex~40_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_19),
	.datad(\rdat1_ex~40_combout ),
	.cin(gnd),
	.combout(rdat1_ex20),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~41 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N28
cycloneive_lcell_comb \rdat1_ex~43 (
// Equation(s):
// rdat1_ex21 = (ccifiwait_0 & (\prif.rdat1_ex [22])) # (!ccifiwait_0 & ((\rdat1_ex~42_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_22),
	.datad(\rdat1_ex~42_combout ),
	.cin(gnd),
	.combout(rdat1_ex21),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~43 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N14
cycloneive_lcell_comb \rdat1_ex~45 (
// Equation(s):
// rdat1_ex22 = (ccifiwait_0 & (\prif.rdat1_ex [21])) # (!ccifiwait_0 & ((\rdat1_ex~44_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_21),
	.datad(\rdat1_ex~44_combout ),
	.cin(gnd),
	.combout(rdat1_ex22),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~45 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N12
cycloneive_lcell_comb \rdat1_ex~47 (
// Equation(s):
// rdat1_ex23 = (ccifiwait_0 & (\prif.rdat1_ex [24])) # (!ccifiwait_0 & ((\rdat1_ex~46_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_24),
	.datad(\rdat1_ex~46_combout ),
	.cin(gnd),
	.combout(rdat1_ex23),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~47 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N2
cycloneive_lcell_comb \rdat1_ex~49 (
// Equation(s):
// rdat1_ex24 = (ccifiwait_0 & (\prif.rdat1_ex [23])) # (!ccifiwait_0 & ((\rdat1_ex~48_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_23),
	.datad(\rdat1_ex~48_combout ),
	.cin(gnd),
	.combout(rdat1_ex24),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~49 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~49 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N0
cycloneive_lcell_comb \rdat1_ex~51 (
// Equation(s):
// rdat1_ex25 = (ccifiwait_0 & (\prif.rdat1_ex [31])) # (!ccifiwait_0 & ((\rdat1_ex~50_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_31),
	.datad(\rdat1_ex~50_combout ),
	.cin(gnd),
	.combout(rdat1_ex25),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~51 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~51 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N26
cycloneive_lcell_comb \rdat1_ex~53 (
// Equation(s):
// rdat1_ex26 = (ccifiwait_0 & (\prif.rdat1_ex [30])) # (!ccifiwait_0 & ((\rdat1_ex~52_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_30),
	.datad(\rdat1_ex~52_combout ),
	.cin(gnd),
	.combout(rdat1_ex26),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~53 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~53 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N24
cycloneive_lcell_comb \rdat1_ex~55 (
// Equation(s):
// rdat1_ex27 = (ccifiwait_0 & (\prif.rdat1_ex [29])) # (!ccifiwait_0 & ((\rdat1_ex~54_combout )))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrdat1_ex_29),
	.datad(\rdat1_ex~54_combout ),
	.cin(gnd),
	.combout(rdat1_ex27),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~55 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~55 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N24
cycloneive_lcell_comb \rdat1_ex~57 (
// Equation(s):
// rdat1_ex28 = (ccifiwait_0 & (\prif.rdat1_ex [26])) # (!ccifiwait_0 & ((\rdat1_ex~56_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_26),
	.datad(\rdat1_ex~56_combout ),
	.cin(gnd),
	.combout(rdat1_ex28),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~57 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~57 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N14
cycloneive_lcell_comb \rdat1_ex~59 (
// Equation(s):
// rdat1_ex29 = (ccifiwait_0 & (\prif.rdat1_ex [25])) # (!ccifiwait_0 & ((\rdat1_ex~58_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_25),
	.datad(\rdat1_ex~58_combout ),
	.cin(gnd),
	.combout(rdat1_ex29),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~59 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~59 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N4
cycloneive_lcell_comb \rdat1_ex~61 (
// Equation(s):
// rdat1_ex30 = (ccifiwait_0 & (\prif.rdat1_ex [28])) # (!ccifiwait_0 & ((\rdat1_ex~60_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_28),
	.datad(\rdat1_ex~60_combout ),
	.cin(gnd),
	.combout(rdat1_ex30),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~61 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~61 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N22
cycloneive_lcell_comb \rdat1_ex~63 (
// Equation(s):
// rdat1_ex31 = (ccifiwait_0 & (\prif.rdat1_ex [27])) # (!ccifiwait_0 & ((\rdat1_ex~62_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrdat1_ex_27),
	.datad(\rdat1_ex~62_combout ),
	.cin(gnd),
	.combout(rdat1_ex31),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~63 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~63 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N10
cycloneive_lcell_comb \ALUScr_ex~13 (
// Equation(s):
// ALUScr_ex2 = (!\prif.imemload_id [28]) # (!Equal15)

	.dataa(gnd),
	.datab(gnd),
	.datac(Equal15),
	.datad(prifimemload_id_28),
	.cin(gnd),
	.combout(ALUScr_ex2),
	.cout());
// synopsys translate_off
defparam \ALUScr_ex~13 .lut_mask = 16'h0FFF;
defparam \ALUScr_ex~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y24_N12
cycloneive_lcell_comb \ALUOP_ex~4 (
// Equation(s):
// ALUOP_ex3 = (!flush_idex & ((ccifiwait_0 & ((\prif.ALUOP_ex [0]))) # (!ccifiwait_0 & (!Selector3))))

	.dataa(flush_idex),
	.datab(Selector3),
	.datac(prifALUOP_ex_0),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(ALUOP_ex3),
	.cout());
// synopsys translate_off
defparam \ALUOP_ex~4 .lut_mask = 16'h5011;
defparam \ALUOP_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N20
cycloneive_lcell_comb \instr_mem~0 (
// Equation(s):
// instr_mem = (exmem_en & ((\prif.instr_ex [3]))) # (!exmem_en & (\prif.instr_mem [3]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_3),
	.datad(prifinstr_ex_3),
	.cin(gnd),
	.combout(instr_mem),
	.cout());
// synopsys translate_off
defparam \instr_mem~0 .lut_mask = 16'hFA50;
defparam \instr_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N6
cycloneive_lcell_comb \instr_mem~1 (
// Equation(s):
// instr_mem1 = (exmem_en & ((\prif.instr_ex [5]))) # (!exmem_en & (\prif.instr_mem [5]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_5),
	.datad(prifinstr_ex_5),
	.cin(gnd),
	.combout(instr_mem1),
	.cout());
// synopsys translate_off
defparam \instr_mem~1 .lut_mask = 16'hFA50;
defparam \instr_mem~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N12
cycloneive_lcell_comb \instr_mem~2 (
// Equation(s):
// instr_mem2 = (exmem_en & ((\prif.instr_ex [4]))) # (!exmem_en & (\prif.instr_mem [4]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifinstr_mem_4),
	.datad(prifinstr_ex_4),
	.cin(gnd),
	.combout(instr_mem2),
	.cout());
// synopsys translate_off
defparam \instr_mem~2 .lut_mask = 16'hFC30;
defparam \instr_mem~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N16
cycloneive_lcell_comb \instr_mem~3 (
// Equation(s):
// instr_mem3 = (exmem_en & ((\prif.instr_ex [2]))) # (!exmem_en & (\prif.instr_mem [2]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_2),
	.datad(prifinstr_ex_2),
	.cin(gnd),
	.combout(instr_mem3),
	.cout());
// synopsys translate_off
defparam \instr_mem~3 .lut_mask = 16'hFA50;
defparam \instr_mem~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N10
cycloneive_lcell_comb \instr_mem~4 (
// Equation(s):
// instr_mem4 = (exmem_en & ((\prif.instr_ex [1]))) # (!exmem_en & (\prif.instr_mem [1]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_1),
	.datad(prifinstr_ex_1),
	.cin(gnd),
	.combout(instr_mem4),
	.cout());
// synopsys translate_off
defparam \instr_mem~4 .lut_mask = 16'hFA50;
defparam \instr_mem~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y30_N28
cycloneive_lcell_comb \instr_mem~5 (
// Equation(s):
// instr_mem5 = (exmem_en & ((\prif.instr_ex [0]))) # (!exmem_en & (\prif.instr_mem [0]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_0),
	.datad(prifinstr_ex_0),
	.cin(gnd),
	.combout(instr_mem5),
	.cout());
// synopsys translate_off
defparam \instr_mem~5 .lut_mask = 16'hFA50;
defparam \instr_mem~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N12
cycloneive_lcell_comb \rdat1_mem~0 (
// Equation(s):
// rdat1_mem = (exmem_en & ((\prif.rdat1_ex [1]))) # (!exmem_en & (\prif.rdat1_mem [1]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifrdat1_mem_1),
	.datad(prifrdat1_ex_1),
	.cin(gnd),
	.combout(rdat1_mem),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~0 .lut_mask = 16'hFA50;
defparam \rdat1_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N30
cycloneive_lcell_comb \PCScr_mem~0 (
// Equation(s):
// PCScr_mem = (exmem_en & (\prif.PCScr_ex [0])) # (!exmem_en & ((\prif.PCScr_mem [0])))

	.dataa(gnd),
	.datab(prifPCScr_ex_0),
	.datac(prifPCScr_mem_0),
	.datad(exmem_en),
	.cin(gnd),
	.combout(PCScr_mem),
	.cout());
// synopsys translate_off
defparam \PCScr_mem~0 .lut_mask = 16'hCCF0;
defparam \PCScr_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N4
cycloneive_lcell_comb \pc_bran_mem~0 (
// Equation(s):
// pc_bran_mem = (exmem_en & ((\prif.pc_ex [1]))) # (!exmem_en & (\prif.pc_bran_mem [1]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifpc_bran_mem_1),
	.datad(prifpc_ex_1),
	.cin(gnd),
	.combout(pc_bran_mem),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~0 .lut_mask = 16'hFA50;
defparam \pc_bran_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N18
cycloneive_lcell_comb \PCScr_mem~1 (
// Equation(s):
// PCScr_mem1 = (exmem_en & ((\prif.PCScr_ex [1]))) # (!exmem_en & (\prif.PCScr_mem [1]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifPCScr_mem_1),
	.datad(prifPCScr_ex_1),
	.cin(gnd),
	.combout(PCScr_mem1),
	.cout());
// synopsys translate_off
defparam \PCScr_mem~1 .lut_mask = 16'hFC30;
defparam \PCScr_mem~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N28
cycloneive_lcell_comb \opcode_ex~0 (
// Equation(s):
// opcode_ex = (ccifiwait_0 & (\prif.opcode_ex [5])) # (!ccifiwait_0 & ((\prif.imemload_id [31])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifopcode_ex_5),
	.datad(prifimemload_id_31),
	.cin(gnd),
	.combout(opcode_ex),
	.cout());
// synopsys translate_off
defparam \opcode_ex~0 .lut_mask = 16'hF3C0;
defparam \opcode_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N4
cycloneive_lcell_comb \opcode_ex~1 (
// Equation(s):
// opcode_ex1 = (ccifiwait_0 & (\prif.opcode_ex [0])) # (!ccifiwait_0 & ((\prif.imemload_id [26])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifopcode_ex_0),
	.datad(prifimemload_id_26),
	.cin(gnd),
	.combout(opcode_ex1),
	.cout());
// synopsys translate_off
defparam \opcode_ex~1 .lut_mask = 16'hF5A0;
defparam \opcode_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N14
cycloneive_lcell_comb \opcode_ex~2 (
// Equation(s):
// opcode_ex2 = (ccifiwait_0 & ((\prif.opcode_ex [1]))) # (!ccifiwait_0 & (\prif.imemload_id [27]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_27),
	.datac(prifopcode_ex_1),
	.datad(gnd),
	.cin(gnd),
	.combout(opcode_ex2),
	.cout());
// synopsys translate_off
defparam \opcode_ex~2 .lut_mask = 16'hE4E4;
defparam \opcode_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N4
cycloneive_lcell_comb \opcode_ex~3 (
// Equation(s):
// opcode_ex3 = (ccifiwait_0 & ((\prif.opcode_ex [2]))) # (!ccifiwait_0 & (\prif.imemload_id [28]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_28),
	.datac(prifopcode_ex_2),
	.datad(gnd),
	.cin(gnd),
	.combout(opcode_ex3),
	.cout());
// synopsys translate_off
defparam \opcode_ex~3 .lut_mask = 16'hE4E4;
defparam \opcode_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N28
cycloneive_lcell_comb \opcode_ex~4 (
// Equation(s):
// opcode_ex4 = (ccifiwait_0 & (\prif.opcode_ex [4])) # (!ccifiwait_0 & ((\prif.imemload_id [30])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifopcode_ex_4),
	.datad(prifimemload_id_30),
	.cin(gnd),
	.combout(opcode_ex4),
	.cout());
// synopsys translate_off
defparam \opcode_ex~4 .lut_mask = 16'hF5A0;
defparam \opcode_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N12
cycloneive_lcell_comb \memren_ex~0 (
// Equation(s):
// memren_ex = (ccifiwait_0 & (((\prif.memren_ex~q )))) # (!ccifiwait_0 & (Equal131 & ((\prif.imemload_id [31]))))

	.dataa(ccifiwait_0),
	.datab(Equal131),
	.datac(prifmemren_ex),
	.datad(prifimemload_id_31),
	.cin(gnd),
	.combout(memren_ex),
	.cout());
// synopsys translate_off
defparam \memren_ex~0 .lut_mask = 16'hE4A0;
defparam \memren_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N26
cycloneive_lcell_comb \memwen_ex~0 (
// Equation(s):
// memwen_ex = (ccifiwait_0 & (\prif.memwen_ex~q )) # (!ccifiwait_0 & ((Equal25)))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifmemwen_ex),
	.datad(Equal25),
	.cin(gnd),
	.combout(memwen_ex),
	.cout());
// synopsys translate_off
defparam \memwen_ex~0 .lut_mask = 16'hF5A0;
defparam \memwen_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N24
cycloneive_lcell_comb \rdat1_mem~1 (
// Equation(s):
// rdat1_mem1 = (exmem_en & ((\prif.rdat1_ex [0]))) # (!exmem_en & (\prif.rdat1_mem [0]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifrdat1_mem_0),
	.datad(prifrdat1_ex_0),
	.cin(gnd),
	.combout(rdat1_mem1),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~1 .lut_mask = 16'hFC30;
defparam \rdat1_mem~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N26
cycloneive_lcell_comb \pc_bran_mem~1 (
// Equation(s):
// pc_bran_mem1 = (exmem_en & ((\prif.pc_ex [0]))) # (!exmem_en & (\prif.pc_bran_mem [0]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_0),
	.datad(prifpc_ex_0),
	.cin(gnd),
	.combout(pc_bran_mem1),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~1 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N12
cycloneive_lcell_comb \rdat1_mem~2 (
// Equation(s):
// rdat1_mem2 = (exmem_en & (\prif.rdat1_ex [3])) # (!exmem_en & ((\prif.rdat1_mem [3])))

	.dataa(prifrdat1_ex_3),
	.datab(gnd),
	.datac(prifrdat1_mem_3),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem2),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~2 .lut_mask = 16'hAAF0;
defparam \rdat1_mem~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N4
cycloneive_lcell_comb \pc_bran_mem~2 (
// Equation(s):
// pc_bran_mem2 = (exmem_en & ((\Add0~2_combout ))) # (!exmem_en & (\prif.pc_bran_mem [3]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_3),
	.datad(Add01),
	.cin(gnd),
	.combout(pc_bran_mem2),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~2 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N14
cycloneive_lcell_comb \rdat1_mem~3 (
// Equation(s):
// rdat1_mem3 = (exmem_en & ((\prif.rdat1_ex [2]))) # (!exmem_en & (\prif.rdat1_mem [2]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifrdat1_mem_2),
	.datad(prifrdat1_ex_2),
	.cin(gnd),
	.combout(rdat1_mem3),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~3 .lut_mask = 16'hFC30;
defparam \rdat1_mem~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N20
cycloneive_lcell_comb \pc_bran_mem~3 (
// Equation(s):
// pc_bran_mem3 = (exmem_en & ((\Add0~0_combout ))) # (!exmem_en & (\prif.pc_bran_mem [2]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_2),
	.datad(Add0),
	.cin(gnd),
	.combout(pc_bran_mem3),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~3 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N20
cycloneive_lcell_comb \rdat1_mem~4 (
// Equation(s):
// rdat1_mem4 = (exmem_en & ((\prif.rdat1_ex [5]))) # (!exmem_en & (\prif.rdat1_mem [5]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifrdat1_mem_5),
	.datad(prifrdat1_ex_5),
	.cin(gnd),
	.combout(rdat1_mem4),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~4 .lut_mask = 16'hFA50;
defparam \rdat1_mem~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N22
cycloneive_lcell_comb \pc_bran_mem~4 (
// Equation(s):
// pc_bran_mem4 = (exmem_en & ((\Add0~6_combout ))) # (!exmem_en & (\prif.pc_bran_mem [5]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_5),
	.datad(Add03),
	.cin(gnd),
	.combout(pc_bran_mem4),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~4 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N8
cycloneive_lcell_comb \rdat1_mem~5 (
// Equation(s):
// rdat1_mem5 = (exmem_en & (\prif.rdat1_ex [4])) # (!exmem_en & ((\prif.rdat1_mem [4])))

	.dataa(prifrdat1_ex_4),
	.datab(exmem_en),
	.datac(prifrdat1_mem_4),
	.datad(gnd),
	.cin(gnd),
	.combout(rdat1_mem5),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~5 .lut_mask = 16'hB8B8;
defparam \rdat1_mem~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y33_N0
cycloneive_lcell_comb \pc_bran_mem~5 (
// Equation(s):
// pc_bran_mem5 = (exmem_en & (\Add0~4_combout )) # (!exmem_en & ((\prif.pc_bran_mem [4])))

	.dataa(Add02),
	.datab(gnd),
	.datac(prifpc_bran_mem_4),
	.datad(exmem_en),
	.cin(gnd),
	.combout(pc_bran_mem5),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~5 .lut_mask = 16'hAAF0;
defparam \pc_bran_mem~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N18
cycloneive_lcell_comb \rdat1_mem~6 (
// Equation(s):
// rdat1_mem6 = (exmem_en & ((\prif.rdat1_ex [7]))) # (!exmem_en & (\prif.rdat1_mem [7]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifrdat1_mem_7),
	.datad(prifrdat1_ex_7),
	.cin(gnd),
	.combout(rdat1_mem6),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~6 .lut_mask = 16'hFC30;
defparam \rdat1_mem~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N30
cycloneive_lcell_comb \pc_bran_mem~6 (
// Equation(s):
// pc_bran_mem6 = (exmem_en & (\Add0~10_combout )) # (!exmem_en & ((\prif.pc_bran_mem [7])))

	.dataa(Add05),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_7),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_bran_mem6),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~6 .lut_mask = 16'hB8B8;
defparam \pc_bran_mem~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N28
cycloneive_lcell_comb \rdat1_mem~7 (
// Equation(s):
// rdat1_mem7 = (exmem_en & (\prif.rdat1_ex [6])) # (!exmem_en & ((\prif.rdat1_mem [6])))

	.dataa(prifrdat1_ex_6),
	.datab(exmem_en),
	.datac(prifrdat1_mem_6),
	.datad(gnd),
	.cin(gnd),
	.combout(rdat1_mem7),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~7 .lut_mask = 16'hB8B8;
defparam \rdat1_mem~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N6
cycloneive_lcell_comb \pc_bran_mem~7 (
// Equation(s):
// pc_bran_mem7 = (exmem_en & ((\Add0~8_combout ))) # (!exmem_en & (\prif.pc_bran_mem [6]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_6),
	.datad(Add04),
	.cin(gnd),
	.combout(pc_bran_mem7),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~7 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N16
cycloneive_lcell_comb \rdat1_mem~8 (
// Equation(s):
// rdat1_mem8 = (exmem_en & (\prif.rdat1_ex [9])) # (!exmem_en & ((\prif.rdat1_mem [9])))

	.dataa(prifrdat1_ex_9),
	.datab(exmem_en),
	.datac(prifrdat1_mem_9),
	.datad(gnd),
	.cin(gnd),
	.combout(rdat1_mem8),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~8 .lut_mask = 16'hB8B8;
defparam \rdat1_mem~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N12
cycloneive_lcell_comb \pc_bran_mem~8 (
// Equation(s):
// pc_bran_mem8 = (exmem_en & ((\Add0~14_combout ))) # (!exmem_en & (\prif.pc_bran_mem [9]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_9),
	.datad(Add07),
	.cin(gnd),
	.combout(pc_bran_mem8),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~8 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N10
cycloneive_lcell_comb \instr_mem~6 (
// Equation(s):
// instr_mem6 = (exmem_en & ((\prif.instr_ex [7]))) # (!exmem_en & (\prif.instr_mem [7]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifinstr_mem_7),
	.datad(prifinstr_ex_7),
	.cin(gnd),
	.combout(instr_mem6),
	.cout());
// synopsys translate_off
defparam \instr_mem~6 .lut_mask = 16'hFC30;
defparam \instr_mem~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N26
cycloneive_lcell_comb \rdat1_mem~9 (
// Equation(s):
// rdat1_mem9 = (exmem_en & ((\prif.rdat1_ex [8]))) # (!exmem_en & (\prif.rdat1_mem [8]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifrdat1_mem_8),
	.datad(prifrdat1_ex_8),
	.cin(gnd),
	.combout(rdat1_mem9),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~9 .lut_mask = 16'hFC30;
defparam \rdat1_mem~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N16
cycloneive_lcell_comb \pc_bran_mem~9 (
// Equation(s):
// pc_bran_mem9 = (exmem_en & ((\Add0~12_combout ))) # (!exmem_en & (\prif.pc_bran_mem [8]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_8),
	.datad(Add06),
	.cin(gnd),
	.combout(pc_bran_mem9),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~9 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N18
cycloneive_lcell_comb \instr_mem~7 (
// Equation(s):
// instr_mem7 = (exmem_en & (\prif.instr_ex [6])) # (!exmem_en & ((\prif.instr_mem [6])))

	.dataa(exmem_en),
	.datab(prifinstr_ex_6),
	.datac(prifinstr_mem_6),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_mem7),
	.cout());
// synopsys translate_off
defparam \instr_mem~7 .lut_mask = 16'hD8D8;
defparam \instr_mem~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N2
cycloneive_lcell_comb \rdat1_mem~10 (
// Equation(s):
// rdat1_mem10 = (exmem_en & ((\prif.rdat1_ex [11]))) # (!exmem_en & (\prif.rdat1_mem [11]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifrdat1_mem_11),
	.datad(prifrdat1_ex_11),
	.cin(gnd),
	.combout(rdat1_mem10),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~10 .lut_mask = 16'hFA50;
defparam \rdat1_mem~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N24
cycloneive_lcell_comb \pc_bran_mem~10 (
// Equation(s):
// pc_bran_mem10 = (exmem_en & ((\Add0~18_combout ))) # (!exmem_en & (\prif.pc_bran_mem [11]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_11),
	.datad(Add09),
	.cin(gnd),
	.combout(pc_bran_mem10),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~10 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N12
cycloneive_lcell_comb \instr_mem~8 (
// Equation(s):
// instr_mem8 = (exmem_en & (\prif.instr_ex [9])) # (!exmem_en & ((\prif.instr_mem [9])))

	.dataa(exmem_en),
	.datab(prifinstr_ex_9),
	.datac(prifinstr_mem_9),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_mem8),
	.cout());
// synopsys translate_off
defparam \instr_mem~8 .lut_mask = 16'hD8D8;
defparam \instr_mem~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N18
cycloneive_lcell_comb \rdat1_mem~11 (
// Equation(s):
// rdat1_mem11 = (exmem_en & (\prif.rdat1_ex [10])) # (!exmem_en & ((\prif.rdat1_mem [10])))

	.dataa(exmem_en),
	.datab(prifrdat1_ex_10),
	.datac(prifrdat1_mem_10),
	.datad(gnd),
	.cin(gnd),
	.combout(rdat1_mem11),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~11 .lut_mask = 16'hD8D8;
defparam \rdat1_mem~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N16
cycloneive_lcell_comb \pc_bran_mem~11 (
// Equation(s):
// pc_bran_mem11 = (exmem_en & ((\Add0~16_combout ))) # (!exmem_en & (\prif.pc_bran_mem [10]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifpc_bran_mem_10),
	.datad(Add08),
	.cin(gnd),
	.combout(pc_bran_mem11),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~11 .lut_mask = 16'hFA50;
defparam \pc_bran_mem~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N6
cycloneive_lcell_comb \instr_mem~9 (
// Equation(s):
// instr_mem9 = (exmem_en & ((\prif.instr_ex [8]))) # (!exmem_en & (\prif.instr_mem [8]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_8),
	.datad(prifinstr_ex_8),
	.cin(gnd),
	.combout(instr_mem9),
	.cout());
// synopsys translate_off
defparam \instr_mem~9 .lut_mask = 16'hFA50;
defparam \instr_mem~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N10
cycloneive_lcell_comb \rdat1_mem~12 (
// Equation(s):
// rdat1_mem12 = (exmem_en & (\prif.rdat1_ex [13])) # (!exmem_en & ((\prif.rdat1_mem [13])))

	.dataa(prifrdat1_ex_13),
	.datab(exmem_en),
	.datac(prifrdat1_mem_13),
	.datad(gnd),
	.cin(gnd),
	.combout(rdat1_mem12),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~12 .lut_mask = 16'hB8B8;
defparam \rdat1_mem~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N24
cycloneive_lcell_comb \pc_bran_mem~12 (
// Equation(s):
// pc_bran_mem12 = (exmem_en & ((\Add0~22_combout ))) # (!exmem_en & (\prif.pc_bran_mem [13]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifpc_bran_mem_13),
	.datad(Add011),
	.cin(gnd),
	.combout(pc_bran_mem12),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~12 .lut_mask = 16'hFA50;
defparam \pc_bran_mem~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N30
cycloneive_lcell_comb \instr_mem~10 (
// Equation(s):
// instr_mem10 = (exmem_en & (\prif.instr_ex [11])) # (!exmem_en & ((\prif.instr_mem [11])))

	.dataa(exmem_en),
	.datab(prifinstr_ex_11),
	.datac(prifinstr_mem_11),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_mem10),
	.cout());
// synopsys translate_off
defparam \instr_mem~10 .lut_mask = 16'hD8D8;
defparam \instr_mem~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N24
cycloneive_lcell_comb \rdat1_mem~13 (
// Equation(s):
// rdat1_mem13 = (exmem_en & ((\prif.rdat1_ex [12]))) # (!exmem_en & (\prif.rdat1_mem [12]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifrdat1_mem_12),
	.datad(prifrdat1_ex_12),
	.cin(gnd),
	.combout(rdat1_mem13),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~13 .lut_mask = 16'hFA50;
defparam \rdat1_mem~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N14
cycloneive_lcell_comb \pc_bran_mem~13 (
// Equation(s):
// pc_bran_mem13 = (exmem_en & ((\Add0~20_combout ))) # (!exmem_en & (\prif.pc_bran_mem [12]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifpc_bran_mem_12),
	.datad(Add010),
	.cin(gnd),
	.combout(pc_bran_mem13),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~13 .lut_mask = 16'hFA50;
defparam \pc_bran_mem~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N0
cycloneive_lcell_comb \instr_mem~11 (
// Equation(s):
// instr_mem11 = (exmem_en & ((\prif.instr_ex [10]))) # (!exmem_en & (\prif.instr_mem [10]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_10),
	.datad(prifinstr_ex_10),
	.cin(gnd),
	.combout(instr_mem11),
	.cout());
// synopsys translate_off
defparam \instr_mem~11 .lut_mask = 16'hFA50;
defparam \instr_mem~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N22
cycloneive_lcell_comb \rdat1_mem~14 (
// Equation(s):
// rdat1_mem14 = (exmem_en & ((\prif.rdat1_ex [15]))) # (!exmem_en & (\prif.rdat1_mem [15]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifrdat1_mem_15),
	.datad(prifrdat1_ex_15),
	.cin(gnd),
	.combout(rdat1_mem14),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~14 .lut_mask = 16'hFA50;
defparam \rdat1_mem~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N6
cycloneive_lcell_comb \pc_bran_mem~14 (
// Equation(s):
// pc_bran_mem14 = (exmem_en & ((\Add0~26_combout ))) # (!exmem_en & (\prif.pc_bran_mem [15]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_15),
	.datad(Add013),
	.cin(gnd),
	.combout(pc_bran_mem14),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~14 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N0
cycloneive_lcell_comb \instr_mem~12 (
// Equation(s):
// instr_mem12 = (exmem_en & ((\prif.instr_ex [13]))) # (!exmem_en & (\prif.instr_mem [13]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_13),
	.datad(prifinstr_ex_13),
	.cin(gnd),
	.combout(instr_mem12),
	.cout());
// synopsys translate_off
defparam \instr_mem~12 .lut_mask = 16'hFA50;
defparam \instr_mem~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N6
cycloneive_lcell_comb \rdat1_mem~15 (
// Equation(s):
// rdat1_mem15 = (exmem_en & ((\prif.rdat1_ex [14]))) # (!exmem_en & (\prif.rdat1_mem [14]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifrdat1_mem_14),
	.datad(prifrdat1_ex_14),
	.cin(gnd),
	.combout(rdat1_mem15),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~15 .lut_mask = 16'hFA50;
defparam \rdat1_mem~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N20
cycloneive_lcell_comb \pc_bran_mem~15 (
// Equation(s):
// pc_bran_mem15 = (exmem_en & ((\Add0~24_combout ))) # (!exmem_en & (\prif.pc_bran_mem [14]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifpc_bran_mem_14),
	.datad(Add012),
	.cin(gnd),
	.combout(pc_bran_mem15),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~15 .lut_mask = 16'hFA50;
defparam \pc_bran_mem~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N2
cycloneive_lcell_comb \instr_mem~13 (
// Equation(s):
// instr_mem13 = (exmem_en & ((\prif.instr_ex [12]))) # (!exmem_en & (\prif.instr_mem [12]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_12),
	.datad(prifinstr_ex_12),
	.cin(gnd),
	.combout(instr_mem13),
	.cout());
// synopsys translate_off
defparam \instr_mem~13 .lut_mask = 16'hFA50;
defparam \instr_mem~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N8
cycloneive_lcell_comb \rdat1_mem~16 (
// Equation(s):
// rdat1_mem16 = (exmem_en & ((\prif.rdat1_ex [23]))) # (!exmem_en & (\prif.rdat1_mem [23]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifrdat1_mem_23),
	.datad(prifrdat1_ex_23),
	.cin(gnd),
	.combout(rdat1_mem16),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~16 .lut_mask = 16'hFA50;
defparam \rdat1_mem~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N30
cycloneive_lcell_comb \pc_bran_mem~16 (
// Equation(s):
// pc_bran_mem16 = (exmem_en & ((\Add0~42_combout ))) # (!exmem_en & (\prif.pc_bran_mem [23]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifpc_bran_mem_23),
	.datad(Add021),
	.cin(gnd),
	.combout(pc_bran_mem16),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~16 .lut_mask = 16'hFA50;
defparam \pc_bran_mem~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N16
cycloneive_lcell_comb \instr_mem~14 (
// Equation(s):
// instr_mem14 = (exmem_en & ((\prif.instr_ex [21]))) # (!exmem_en & (\prif.instr_mem [21]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_21),
	.datad(prifinstr_ex_21),
	.cin(gnd),
	.combout(instr_mem14),
	.cout());
// synopsys translate_off
defparam \instr_mem~14 .lut_mask = 16'hFA50;
defparam \instr_mem~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N20
cycloneive_lcell_comb \rdat1_mem~17 (
// Equation(s):
// rdat1_mem17 = (exmem_en & (\prif.rdat1_ex [22])) # (!exmem_en & ((\prif.rdat1_mem [22])))

	.dataa(gnd),
	.datab(prifrdat1_ex_22),
	.datac(prifrdat1_mem_22),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem17),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~17 .lut_mask = 16'hCCF0;
defparam \rdat1_mem~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N10
cycloneive_lcell_comb \pc_bran_mem~17 (
// Equation(s):
// pc_bran_mem17 = (exmem_en & ((\Add0~40_combout ))) # (!exmem_en & (\prif.pc_bran_mem [22]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_22),
	.datad(Add020),
	.cin(gnd),
	.combout(pc_bran_mem17),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~17 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y28_N8
cycloneive_lcell_comb \instr_mem~15 (
// Equation(s):
// instr_mem15 = (exmem_en & ((\prif.instr_ex [20]))) # (!exmem_en & (\prif.instr_mem [20]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_20),
	.datad(prifinstr_ex_20),
	.cin(gnd),
	.combout(instr_mem15),
	.cout());
// synopsys translate_off
defparam \instr_mem~15 .lut_mask = 16'hFA50;
defparam \instr_mem~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N16
cycloneive_lcell_comb \rdat1_mem~18 (
// Equation(s):
// rdat1_mem18 = (exmem_en & (\prif.rdat1_ex [21])) # (!exmem_en & ((\prif.rdat1_mem [21])))

	.dataa(gnd),
	.datab(prifrdat1_ex_21),
	.datac(prifrdat1_mem_21),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem18),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~18 .lut_mask = 16'hCCF0;
defparam \rdat1_mem~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N18
cycloneive_lcell_comb \pc_bran_mem~18 (
// Equation(s):
// pc_bran_mem18 = (exmem_en & (\Add0~38_combout )) # (!exmem_en & ((\prif.pc_bran_mem [21])))

	.dataa(gnd),
	.datab(Add019),
	.datac(prifpc_bran_mem_21),
	.datad(exmem_en),
	.cin(gnd),
	.combout(pc_bran_mem18),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~18 .lut_mask = 16'hCCF0;
defparam \pc_bran_mem~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N0
cycloneive_lcell_comb \instr_mem~16 (
// Equation(s):
// instr_mem16 = (exmem_en & (\prif.instr_ex [19])) # (!exmem_en & ((\prif.instr_mem [19])))

	.dataa(prifinstr_ex_19),
	.datab(gnd),
	.datac(prifinstr_mem_19),
	.datad(exmem_en),
	.cin(gnd),
	.combout(instr_mem16),
	.cout());
// synopsys translate_off
defparam \instr_mem~16 .lut_mask = 16'hAAF0;
defparam \instr_mem~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N24
cycloneive_lcell_comb \rdat1_mem~19 (
// Equation(s):
// rdat1_mem19 = (exmem_en & ((\prif.rdat1_ex [29]))) # (!exmem_en & (\prif.rdat1_mem [29]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifrdat1_mem_29),
	.datad(prifrdat1_ex_29),
	.cin(gnd),
	.combout(rdat1_mem19),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~19 .lut_mask = 16'hFA50;
defparam \rdat1_mem~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y32_N30
cycloneive_lcell_comb \pc_bran_mem~19 (
// Equation(s):
// pc_bran_mem19 = (exmem_en & ((\Add0~54_combout ))) # (!exmem_en & (\prif.pc_bran_mem [29]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifpc_bran_mem_29),
	.datad(Add027),
	.cin(gnd),
	.combout(pc_bran_mem19),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~19 .lut_mask = 16'hFA50;
defparam \pc_bran_mem~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y31_N6
cycloneive_lcell_comb \prif.pc_mem[29]~0 (
// Equation(s):
// prifpc_mem_291 = (\prif.pc_mem[15]~0_combout  & ((\prif.pc_mem [29]))) # (!\prif.pc_mem[15]~0_combout  & (\prif.pc_ex [29]))

	.dataa(prifpc_ex_29),
	.datab(gnd),
	.datac(prifpc_mem_29),
	.datad(prifpc_mem_151),
	.cin(gnd),
	.combout(prifpc_mem_291),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[29]~0 .lut_mask = 16'hF0AA;
defparam \prif.pc_mem[29]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N2
cycloneive_lcell_comb \rdat1_mem~20 (
// Equation(s):
// rdat1_mem20 = (exmem_en & (\prif.rdat1_ex [28])) # (!exmem_en & ((\prif.rdat1_mem [28])))

	.dataa(gnd),
	.datab(prifrdat1_ex_28),
	.datac(prifrdat1_mem_28),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem20),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~20 .lut_mask = 16'hCCF0;
defparam \rdat1_mem~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N4
cycloneive_lcell_comb \pc_bran_mem~20 (
// Equation(s):
// pc_bran_mem20 = (exmem_en & (\Add0~52_combout )) # (!exmem_en & ((\prif.pc_bran_mem [28])))

	.dataa(gnd),
	.datab(Add026),
	.datac(prifpc_bran_mem_28),
	.datad(exmem_en),
	.cin(gnd),
	.combout(pc_bran_mem20),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~20 .lut_mask = 16'hCCF0;
defparam \pc_bran_mem~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N4
cycloneive_lcell_comb \prif.pc_mem[28]~1 (
// Equation(s):
// prifpc_mem_281 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [28])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [28])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_28),
	.datad(prifpc_ex_28),
	.cin(gnd),
	.combout(prifpc_mem_281),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[28]~1 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[28]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N14
cycloneive_lcell_comb \rdat1_mem~21 (
// Equation(s):
// rdat1_mem21 = (exmem_en & (\prif.rdat1_ex [31])) # (!exmem_en & ((\prif.rdat1_mem [31])))

	.dataa(prifrdat1_ex_31),
	.datab(gnd),
	.datac(prifrdat1_mem_31),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem21),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~21 .lut_mask = 16'hAAF0;
defparam \rdat1_mem~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N12
cycloneive_lcell_comb \pc_bran_mem~21 (
// Equation(s):
// pc_bran_mem21 = (exmem_en & (\Add0~58_combout )) # (!exmem_en & ((\prif.pc_bran_mem [31])))

	.dataa(gnd),
	.datab(Add029),
	.datac(prifpc_bran_mem_31),
	.datad(exmem_en),
	.cin(gnd),
	.combout(pc_bran_mem21),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~21 .lut_mask = 16'hCCF0;
defparam \pc_bran_mem~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N22
cycloneive_lcell_comb \prif.pc_mem[31]~2 (
// Equation(s):
// prifpc_mem_311 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [31])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [31])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_31),
	.datad(prifpc_ex_31),
	.cin(gnd),
	.combout(prifpc_mem_311),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[31]~2 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[31]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y33_N30
cycloneive_lcell_comb \rdat1_mem~22 (
// Equation(s):
// rdat1_mem22 = (exmem_en & (\prif.rdat1_ex [30])) # (!exmem_en & ((\prif.rdat1_mem [30])))

	.dataa(prifrdat1_ex_30),
	.datab(gnd),
	.datac(prifrdat1_mem_30),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem22),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~22 .lut_mask = 16'hAAF0;
defparam \rdat1_mem~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N24
cycloneive_lcell_comb \pc_bran_mem~22 (
// Equation(s):
// pc_bran_mem22 = (exmem_en & (\Add0~56_combout )) # (!exmem_en & ((\prif.pc_bran_mem [30])))

	.dataa(Add028),
	.datab(gnd),
	.datac(prifpc_bran_mem_30),
	.datad(exmem_en),
	.cin(gnd),
	.combout(pc_bran_mem22),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~22 .lut_mask = 16'hAAF0;
defparam \pc_bran_mem~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N24
cycloneive_lcell_comb \prif.pc_mem[30]~3 (
// Equation(s):
// prifpc_mem_301 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [30])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [30])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_30),
	.datad(prifpc_ex_30),
	.cin(gnd),
	.combout(prifpc_mem_301),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[30]~3 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[30]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N20
cycloneive_lcell_comb \rdat1_mem~23 (
// Equation(s):
// rdat1_mem23 = (exmem_en & (\prif.rdat1_ex [20])) # (!exmem_en & ((\prif.rdat1_mem [20])))

	.dataa(gnd),
	.datab(prifrdat1_ex_20),
	.datac(prifrdat1_mem_20),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem23),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~23 .lut_mask = 16'hCCF0;
defparam \rdat1_mem~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N22
cycloneive_lcell_comb \pc_bran_mem~23 (
// Equation(s):
// pc_bran_mem23 = (exmem_en & ((\Add0~36_combout ))) # (!exmem_en & (\prif.pc_bran_mem [20]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_20),
	.datad(Add018),
	.cin(gnd),
	.combout(pc_bran_mem23),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~23 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N16
cycloneive_lcell_comb \instr_mem~17 (
// Equation(s):
// instr_mem17 = (exmem_en & ((\prif.instr_ex [18]))) # (!exmem_en & (\prif.instr_mem [18]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifinstr_mem_18),
	.datad(prifinstr_ex_18),
	.cin(gnd),
	.combout(instr_mem17),
	.cout());
// synopsys translate_off
defparam \instr_mem~17 .lut_mask = 16'hFC30;
defparam \instr_mem~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N4
cycloneive_lcell_comb \rdat1_mem~24 (
// Equation(s):
// rdat1_mem24 = (exmem_en & (\prif.rdat1_ex [17])) # (!exmem_en & ((\prif.rdat1_mem [17])))

	.dataa(gnd),
	.datab(prifrdat1_ex_17),
	.datac(prifrdat1_mem_17),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem24),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~24 .lut_mask = 16'hCCF0;
defparam \rdat1_mem~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N2
cycloneive_lcell_comb \pc_bran_mem~24 (
// Equation(s):
// pc_bran_mem24 = (exmem_en & ((\Add0~30_combout ))) # (!exmem_en & (\prif.pc_bran_mem [17]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_17),
	.datad(Add015),
	.cin(gnd),
	.combout(pc_bran_mem24),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~24 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N8
cycloneive_lcell_comb \instr_mem~18 (
// Equation(s):
// instr_mem18 = (exmem_en & ((\prif.instr_ex [15]))) # (!exmem_en & (\prif.instr_mem [15]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifinstr_mem_15),
	.datad(prifinstr_ex_15),
	.cin(gnd),
	.combout(instr_mem18),
	.cout());
// synopsys translate_off
defparam \instr_mem~18 .lut_mask = 16'hFC30;
defparam \instr_mem~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N14
cycloneive_lcell_comb \rdat1_mem~25 (
// Equation(s):
// rdat1_mem25 = (exmem_en & ((\prif.rdat1_ex [16]))) # (!exmem_en & (\prif.rdat1_mem [16]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifrdat1_mem_16),
	.datad(prifrdat1_ex_16),
	.cin(gnd),
	.combout(rdat1_mem25),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~25 .lut_mask = 16'hFC30;
defparam \rdat1_mem~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N28
cycloneive_lcell_comb \pc_bran_mem~25 (
// Equation(s):
// pc_bran_mem25 = (exmem_en & ((\Add0~28_combout ))) # (!exmem_en & (\prif.pc_bran_mem [16]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_16),
	.datad(Add014),
	.cin(gnd),
	.combout(pc_bran_mem25),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~25 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y31_N26
cycloneive_lcell_comb \instr_mem~19 (
// Equation(s):
// instr_mem19 = (exmem_en & (\prif.instr_ex [14])) # (!exmem_en & ((\prif.instr_mem [14])))

	.dataa(prifinstr_ex_14),
	.datab(exmem_en),
	.datac(prifinstr_mem_14),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_mem19),
	.cout());
// synopsys translate_off
defparam \instr_mem~19 .lut_mask = 16'hB8B8;
defparam \instr_mem~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N10
cycloneive_lcell_comb \rdat1_mem~26 (
// Equation(s):
// rdat1_mem26 = (exmem_en & (\prif.rdat1_ex [19])) # (!exmem_en & ((\prif.rdat1_mem [19])))

	.dataa(prifrdat1_ex_19),
	.datab(gnd),
	.datac(prifrdat1_mem_19),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem26),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~26 .lut_mask = 16'hAAF0;
defparam \rdat1_mem~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N18
cycloneive_lcell_comb \pc_bran_mem~26 (
// Equation(s):
// pc_bran_mem26 = (exmem_en & ((\Add0~34_combout ))) # (!exmem_en & (\prif.pc_bran_mem [19]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_19),
	.datad(Add017),
	.cin(gnd),
	.combout(pc_bran_mem26),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~26 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N0
cycloneive_lcell_comb \instr_mem~20 (
// Equation(s):
// instr_mem20 = (exmem_en & (\prif.instr_ex [17])) # (!exmem_en & ((\prif.instr_mem [17])))

	.dataa(exmem_en),
	.datab(prifinstr_ex_17),
	.datac(prifinstr_mem_17),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_mem20),
	.cout());
// synopsys translate_off
defparam \instr_mem~20 .lut_mask = 16'hD8D8;
defparam \instr_mem~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N2
cycloneive_lcell_comb \rdat1_mem~27 (
// Equation(s):
// rdat1_mem27 = (exmem_en & ((\prif.rdat1_ex [18]))) # (!exmem_en & (\prif.rdat1_mem [18]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifrdat1_mem_18),
	.datad(prifrdat1_ex_18),
	.cin(gnd),
	.combout(rdat1_mem27),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~27 .lut_mask = 16'hFA50;
defparam \rdat1_mem~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N8
cycloneive_lcell_comb \pc_bran_mem~27 (
// Equation(s):
// pc_bran_mem27 = (exmem_en & ((\Add0~32_combout ))) # (!exmem_en & (\prif.pc_bran_mem [18]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifpc_bran_mem_18),
	.datad(Add016),
	.cin(gnd),
	.combout(pc_bran_mem27),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~27 .lut_mask = 16'hFA50;
defparam \pc_bran_mem~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N10
cycloneive_lcell_comb \instr_mem~21 (
// Equation(s):
// instr_mem21 = (exmem_en & ((\prif.instr_ex [16]))) # (!exmem_en & (\prif.instr_mem [16]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifinstr_mem_16),
	.datad(prifinstr_ex_16),
	.cin(gnd),
	.combout(instr_mem21),
	.cout());
// synopsys translate_off
defparam \instr_mem~21 .lut_mask = 16'hFA50;
defparam \instr_mem~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N0
cycloneive_lcell_comb \rdat1_mem~28 (
// Equation(s):
// rdat1_mem28 = (exmem_en & ((\prif.rdat1_ex [25]))) # (!exmem_en & (\prif.rdat1_mem [25]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifrdat1_mem_25),
	.datad(prifrdat1_ex_25),
	.cin(gnd),
	.combout(rdat1_mem28),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~28 .lut_mask = 16'hFC30;
defparam \rdat1_mem~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N26
cycloneive_lcell_comb \pc_bran_mem~28 (
// Equation(s):
// pc_bran_mem28 = (exmem_en & ((\Add0~46_combout ))) # (!exmem_en & (\prif.pc_bran_mem [25]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_25),
	.datad(Add023),
	.cin(gnd),
	.combout(pc_bran_mem28),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~28 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N12
cycloneive_lcell_comb \instr_mem~22 (
// Equation(s):
// instr_mem22 = (exmem_en & ((\prif.instr_ex [23]))) # (!exmem_en & (\prif.instr_mem [23]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifinstr_mem_23),
	.datad(prifinstr_ex_23),
	.cin(gnd),
	.combout(instr_mem22),
	.cout());
// synopsys translate_off
defparam \instr_mem~22 .lut_mask = 16'hFC30;
defparam \instr_mem~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N2
cycloneive_lcell_comb \rdat1_mem~29 (
// Equation(s):
// rdat1_mem29 = (exmem_en & (\prif.rdat1_ex [24])) # (!exmem_en & ((\prif.rdat1_mem [24])))

	.dataa(gnd),
	.datab(prifrdat1_ex_24),
	.datac(prifrdat1_mem_24),
	.datad(exmem_en),
	.cin(gnd),
	.combout(rdat1_mem29),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~29 .lut_mask = 16'hCCF0;
defparam \rdat1_mem~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N28
cycloneive_lcell_comb \pc_bran_mem~29 (
// Equation(s):
// pc_bran_mem29 = (exmem_en & ((\Add0~44_combout ))) # (!exmem_en & (\prif.pc_bran_mem [24]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_24),
	.datad(Add022),
	.cin(gnd),
	.combout(pc_bran_mem29),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~29 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N14
cycloneive_lcell_comb \instr_mem~23 (
// Equation(s):
// instr_mem23 = (exmem_en & ((\prif.instr_ex [22]))) # (!exmem_en & (\prif.instr_mem [22]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifinstr_mem_22),
	.datad(prifinstr_ex_22),
	.cin(gnd),
	.combout(instr_mem23),
	.cout());
// synopsys translate_off
defparam \instr_mem~23 .lut_mask = 16'hFC30;
defparam \instr_mem~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N6
cycloneive_lcell_comb \rdat1_mem~30 (
// Equation(s):
// rdat1_mem30 = (exmem_en & ((\prif.rdat1_ex [27]))) # (!exmem_en & (\prif.rdat1_mem [27]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifrdat1_mem_27),
	.datad(prifrdat1_ex_27),
	.cin(gnd),
	.combout(rdat1_mem30),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~30 .lut_mask = 16'hFC30;
defparam \rdat1_mem~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N16
cycloneive_lcell_comb \pc_bran_mem~30 (
// Equation(s):
// pc_bran_mem30 = (exmem_en & ((\Add0~50_combout ))) # (!exmem_en & (\prif.pc_bran_mem [27]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifpc_bran_mem_27),
	.datad(Add025),
	.cin(gnd),
	.combout(pc_bran_mem30),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~30 .lut_mask = 16'hFC30;
defparam \pc_bran_mem~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y32_N30
cycloneive_lcell_comb \instr_mem~24 (
// Equation(s):
// instr_mem24 = (exmem_en & ((\prif.instr_ex [25]))) # (!exmem_en & (\prif.instr_mem [25]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifinstr_mem_25),
	.datad(prifinstr_ex_25),
	.cin(gnd),
	.combout(instr_mem24),
	.cout());
// synopsys translate_off
defparam \instr_mem~24 .lut_mask = 16'hFC30;
defparam \instr_mem~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N28
cycloneive_lcell_comb \rdat1_mem~31 (
// Equation(s):
// rdat1_mem31 = (exmem_en & (\prif.rdat1_ex [26])) # (!exmem_en & ((\prif.rdat1_mem [26])))

	.dataa(exmem_en),
	.datab(prifrdat1_ex_26),
	.datac(prifrdat1_mem_26),
	.datad(gnd),
	.cin(gnd),
	.combout(rdat1_mem31),
	.cout());
// synopsys translate_off
defparam \rdat1_mem~31 .lut_mask = 16'hD8D8;
defparam \rdat1_mem~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N14
cycloneive_lcell_comb \pc_bran_mem~31 (
// Equation(s):
// pc_bran_mem31 = (exmem_en & ((\Add0~48_combout ))) # (!exmem_en & (\prif.pc_bran_mem [26]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifpc_bran_mem_26),
	.datad(Add024),
	.cin(gnd),
	.combout(pc_bran_mem31),
	.cout());
// synopsys translate_off
defparam \pc_bran_mem~31 .lut_mask = 16'hFA50;
defparam \pc_bran_mem~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y32_N24
cycloneive_lcell_comb \instr_mem~25 (
// Equation(s):
// instr_mem25 = (exmem_en & (\prif.instr_ex [24])) # (!exmem_en & ((\prif.instr_mem [24])))

	.dataa(exmem_en),
	.datab(prifinstr_ex_24),
	.datac(prifinstr_mem_24),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_mem25),
	.cout());
// synopsys translate_off
defparam \instr_mem~25 .lut_mask = 16'hD8D8;
defparam \instr_mem~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N18
cycloneive_lcell_comb \dmemstore~1 (
// Equation(s):
// dmemstore1 = (exmem_en & ((\Mux62~0_combout ) # ((\Mux62~1_combout )))) # (!exmem_en & (((prifdmemstore_1))))

	.dataa(exmem_en),
	.datab(Mux62),
	.datac(prifdmemstore_1),
	.datad(Mux621),
	.cin(gnd),
	.combout(dmemstore1),
	.cout());
// synopsys translate_off
defparam \dmemstore~1 .lut_mask = 16'hFAD8;
defparam \dmemstore~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N20
cycloneive_lcell_comb \dmemstore~2 (
// Equation(s):
// dmemstore2 = (exmem_en & ((\Mux61~1_combout ))) # (!exmem_en & (prifdmemstore_2))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_2),
	.datad(Mux61),
	.cin(gnd),
	.combout(dmemstore2),
	.cout());
// synopsys translate_off
defparam \dmemstore~2 .lut_mask = 16'hFA50;
defparam \dmemstore~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N26
cycloneive_lcell_comb \dmemstore~3 (
// Equation(s):
// dmemstore3 = (exmem_en & ((\Mux60~1_combout ))) # (!exmem_en & (prifdmemstore_3))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_3),
	.datad(Mux602),
	.cin(gnd),
	.combout(dmemstore3),
	.cout());
// synopsys translate_off
defparam \dmemstore~3 .lut_mask = 16'hFA50;
defparam \dmemstore~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N16
cycloneive_lcell_comb \dmemstore~4 (
// Equation(s):
// dmemstore4 = (exmem_en & (\Mux59~1_combout )) # (!exmem_en & ((prifdmemstore_4)))

	.dataa(exmem_en),
	.datab(Mux592),
	.datac(prifdmemstore_4),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemstore4),
	.cout());
// synopsys translate_off
defparam \dmemstore~4 .lut_mask = 16'hD8D8;
defparam \dmemstore~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N2
cycloneive_lcell_comb \dmemstore~5 (
// Equation(s):
// dmemstore5 = (exmem_en & ((\Mux58~1_combout ))) # (!exmem_en & (prifdmemstore_5))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_5),
	.datad(Mux582),
	.cin(gnd),
	.combout(dmemstore5),
	.cout());
// synopsys translate_off
defparam \dmemstore~5 .lut_mask = 16'hFA50;
defparam \dmemstore~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N24
cycloneive_lcell_comb \dmemstore~6 (
// Equation(s):
// dmemstore6 = (exmem_en & ((\Mux57~1_combout ))) # (!exmem_en & (prifdmemstore_6))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_6),
	.datad(Mux572),
	.cin(gnd),
	.combout(dmemstore6),
	.cout());
// synopsys translate_off
defparam \dmemstore~6 .lut_mask = 16'hFA50;
defparam \dmemstore~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N20
cycloneive_lcell_comb \dmemstore~7 (
// Equation(s):
// dmemstore7 = (exmem_en & (\Mux56~1_combout )) # (!exmem_en & ((prifdmemstore_7)))

	.dataa(Mux562),
	.datab(exmem_en),
	.datac(prifdmemstore_7),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemstore7),
	.cout());
// synopsys translate_off
defparam \dmemstore~7 .lut_mask = 16'hB8B8;
defparam \dmemstore~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N10
cycloneive_lcell_comb \dmemstore~8 (
// Equation(s):
// dmemstore8 = (exmem_en & (\Mux55~1_combout )) # (!exmem_en & ((prifdmemstore_8)))

	.dataa(exmem_en),
	.datab(Mux552),
	.datac(prifdmemstore_8),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemstore8),
	.cout());
// synopsys translate_off
defparam \dmemstore~8 .lut_mask = 16'hD8D8;
defparam \dmemstore~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N18
cycloneive_lcell_comb \dmemstore~9 (
// Equation(s):
// dmemstore9 = (exmem_en & ((\Mux54~1_combout ))) # (!exmem_en & (prifdmemstore_9))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemstore_9),
	.datad(Mux542),
	.cin(gnd),
	.combout(dmemstore9),
	.cout());
// synopsys translate_off
defparam \dmemstore~9 .lut_mask = 16'hFC30;
defparam \dmemstore~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N20
cycloneive_lcell_comb \dmemstore~10 (
// Equation(s):
// dmemstore10 = (exmem_en & ((\Mux53~1_combout ))) # (!exmem_en & (prifdmemstore_10))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_10),
	.datad(Mux532),
	.cin(gnd),
	.combout(dmemstore10),
	.cout());
// synopsys translate_off
defparam \dmemstore~10 .lut_mask = 16'hFA50;
defparam \dmemstore~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N6
cycloneive_lcell_comb \dmemstore~11 (
// Equation(s):
// dmemstore11 = (exmem_en & (\Mux52~1_combout )) # (!exmem_en & ((prifdmemstore_11)))

	.dataa(exmem_en),
	.datab(Mux522),
	.datac(prifdmemstore_11),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemstore11),
	.cout());
// synopsys translate_off
defparam \dmemstore~11 .lut_mask = 16'hD8D8;
defparam \dmemstore~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N28
cycloneive_lcell_comb \dmemstore~12 (
// Equation(s):
// dmemstore12 = (exmem_en & ((\Mux51~1_combout ))) # (!exmem_en & (prifdmemstore_12))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_12),
	.datad(Mux512),
	.cin(gnd),
	.combout(dmemstore12),
	.cout());
// synopsys translate_off
defparam \dmemstore~12 .lut_mask = 16'hFA50;
defparam \dmemstore~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y26_N12
cycloneive_lcell_comb \dmemstore~13 (
// Equation(s):
// dmemstore13 = (exmem_en & ((\Mux50~1_combout ))) # (!exmem_en & (prifdmemstore_13))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_13),
	.datad(Mux502),
	.cin(gnd),
	.combout(dmemstore13),
	.cout());
// synopsys translate_off
defparam \dmemstore~13 .lut_mask = 16'hFA50;
defparam \dmemstore~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N18
cycloneive_lcell_comb \dmemstore~14 (
// Equation(s):
// dmemstore14 = (exmem_en & ((\Mux49~1_combout ))) # (!exmem_en & (prifdmemstore_14))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_14),
	.datad(Mux492),
	.cin(gnd),
	.combout(dmemstore14),
	.cout());
// synopsys translate_off
defparam \dmemstore~14 .lut_mask = 16'hFA50;
defparam \dmemstore~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N24
cycloneive_lcell_comb \dmemstore~15 (
// Equation(s):
// dmemstore15 = (exmem_en & (\Mux48~1_combout )) # (!exmem_en & ((prifdmemstore_15)))

	.dataa(exmem_en),
	.datab(Mux482),
	.datac(prifdmemstore_15),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemstore15),
	.cout());
// synopsys translate_off
defparam \dmemstore~15 .lut_mask = 16'hD8D8;
defparam \dmemstore~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N10
cycloneive_lcell_comb \dmemstore~16 (
// Equation(s):
// dmemstore16 = (exmem_en & ((\Mux47~1_combout ))) # (!exmem_en & (prifdmemstore_16))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_16),
	.datad(Mux47),
	.cin(gnd),
	.combout(dmemstore16),
	.cout());
// synopsys translate_off
defparam \dmemstore~16 .lut_mask = 16'hFA50;
defparam \dmemstore~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N12
cycloneive_lcell_comb \dmemstore~17 (
// Equation(s):
// dmemstore17 = (exmem_en & ((\Mux46~1_combout ))) # (!exmem_en & (prifdmemstore_17))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_17),
	.datad(Mux46),
	.cin(gnd),
	.combout(dmemstore17),
	.cout());
// synopsys translate_off
defparam \dmemstore~17 .lut_mask = 16'hFA50;
defparam \dmemstore~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y30_N2
cycloneive_lcell_comb \dmemstore~18 (
// Equation(s):
// dmemstore18 = (exmem_en & ((\Mux45~1_combout ))) # (!exmem_en & (prifdmemstore_18))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_18),
	.datad(Mux45),
	.cin(gnd),
	.combout(dmemstore18),
	.cout());
// synopsys translate_off
defparam \dmemstore~18 .lut_mask = 16'hFA50;
defparam \dmemstore~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N20
cycloneive_lcell_comb \dmemstore~19 (
// Equation(s):
// dmemstore19 = (exmem_en & ((\Mux44~1_combout ))) # (!exmem_en & (prifdmemstore_19))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemstore_19),
	.datad(Mux44),
	.cin(gnd),
	.combout(dmemstore19),
	.cout());
// synopsys translate_off
defparam \dmemstore~19 .lut_mask = 16'hFC30;
defparam \dmemstore~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N6
cycloneive_lcell_comb \dmemstore~20 (
// Equation(s):
// dmemstore20 = (exmem_en & (\Mux43~1_combout )) # (!exmem_en & ((prifdmemstore_20)))

	.dataa(Mux43),
	.datab(gnd),
	.datac(prifdmemstore_20),
	.datad(exmem_en),
	.cin(gnd),
	.combout(dmemstore20),
	.cout());
// synopsys translate_off
defparam \dmemstore~20 .lut_mask = 16'hAAF0;
defparam \dmemstore~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N12
cycloneive_lcell_comb \dmemstore~21 (
// Equation(s):
// dmemstore21 = (exmem_en & ((\Mux42~1_combout ))) # (!exmem_en & (prifdmemstore_21))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemstore_21),
	.datad(Mux42),
	.cin(gnd),
	.combout(dmemstore21),
	.cout());
// synopsys translate_off
defparam \dmemstore~21 .lut_mask = 16'hFC30;
defparam \dmemstore~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N30
cycloneive_lcell_comb \dmemstore~22 (
// Equation(s):
// dmemstore22 = (exmem_en & ((\Mux41~1_combout ))) # (!exmem_en & (prifdmemstore_22))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemstore_22),
	.datad(Mux41),
	.cin(gnd),
	.combout(dmemstore22),
	.cout());
// synopsys translate_off
defparam \dmemstore~22 .lut_mask = 16'hFC30;
defparam \dmemstore~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N10
cycloneive_lcell_comb \dmemstore~23 (
// Equation(s):
// dmemstore23 = (exmem_en & (\Mux40~1_combout )) # (!exmem_en & ((prifdmemstore_23)))

	.dataa(Mux40),
	.datab(exmem_en),
	.datac(prifdmemstore_23),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemstore23),
	.cout());
// synopsys translate_off
defparam \dmemstore~23 .lut_mask = 16'hB8B8;
defparam \dmemstore~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y27_N0
cycloneive_lcell_comb \dmemstore~24 (
// Equation(s):
// dmemstore24 = (exmem_en & ((\Mux39~1_combout ))) # (!exmem_en & (prifdmemstore_24))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_24),
	.datad(Mux39),
	.cin(gnd),
	.combout(dmemstore24),
	.cout());
// synopsys translate_off
defparam \dmemstore~24 .lut_mask = 16'hFA50;
defparam \dmemstore~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N16
cycloneive_lcell_comb \dmemstore~25 (
// Equation(s):
// dmemstore25 = (exmem_en & ((\Mux38~1_combout ))) # (!exmem_en & (prifdmemstore_25))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemstore_25),
	.datad(Mux38),
	.cin(gnd),
	.combout(dmemstore25),
	.cout());
// synopsys translate_off
defparam \dmemstore~25 .lut_mask = 16'hFC30;
defparam \dmemstore~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y27_N2
cycloneive_lcell_comb \dmemstore~26 (
// Equation(s):
// dmemstore26 = (exmem_en & ((\Mux37~1_combout ))) # (!exmem_en & (prifdmemstore_26))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemstore_26),
	.datad(Mux37),
	.cin(gnd),
	.combout(dmemstore26),
	.cout());
// synopsys translate_off
defparam \dmemstore~26 .lut_mask = 16'hFC30;
defparam \dmemstore~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y26_N26
cycloneive_lcell_comb \dmemstore~27 (
// Equation(s):
// dmemstore27 = (exmem_en & ((\Mux36~1_combout ))) # (!exmem_en & (prifdmemstore_27))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemstore_27),
	.datad(Mux36),
	.cin(gnd),
	.combout(dmemstore27),
	.cout());
// synopsys translate_off
defparam \dmemstore~27 .lut_mask = 16'hFC30;
defparam \dmemstore~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y26_N18
cycloneive_lcell_comb \dmemstore~28 (
// Equation(s):
// dmemstore28 = (exmem_en & ((\Mux35~1_combout ))) # (!exmem_en & (prifdmemstore_28))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdmemstore_28),
	.datad(Mux35),
	.cin(gnd),
	.combout(dmemstore28),
	.cout());
// synopsys translate_off
defparam \dmemstore~28 .lut_mask = 16'hFA50;
defparam \dmemstore~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y30_N2
cycloneive_lcell_comb \dmemstore~29 (
// Equation(s):
// dmemstore29 = (exmem_en & ((\Mux34~1_combout ))) # (!exmem_en & (prifdmemstore_29))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemstore_29),
	.datad(Mux34),
	.cin(gnd),
	.combout(dmemstore29),
	.cout());
// synopsys translate_off
defparam \dmemstore~29 .lut_mask = 16'hFC30;
defparam \dmemstore~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y28_N22
cycloneive_lcell_comb \dmemstore~30 (
// Equation(s):
// dmemstore30 = (exmem_en & (\Mux33~1_combout )) # (!exmem_en & ((prifdmemstore_30)))

	.dataa(exmem_en),
	.datab(Mux33),
	.datac(prifdmemstore_30),
	.datad(gnd),
	.cin(gnd),
	.combout(dmemstore30),
	.cout());
// synopsys translate_off
defparam \dmemstore~30 .lut_mask = 16'hD8D8;
defparam \dmemstore~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N8
cycloneive_lcell_comb \dmemstore~31 (
// Equation(s):
// dmemstore31 = (exmem_en & ((\Mux32~1_combout ))) # (!exmem_en & (prifdmemstore_31))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdmemstore_31),
	.datad(Mux32),
	.cin(gnd),
	.combout(dmemstore31),
	.cout());
// synopsys translate_off
defparam \dmemstore~31 .lut_mask = 16'hFC30;
defparam \dmemstore~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N14
cycloneive_lcell_comb \halt_ex~0 (
// Equation(s):
// halt_ex = (ccifiwait_0 & ((\prif.halt_ex~q ))) # (!ccifiwait_0 & (Equal26))

	.dataa(Equal26),
	.datab(gnd),
	.datac(prifhalt_ex),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(halt_ex),
	.cout());
// synopsys translate_off
defparam \halt_ex~0 .lut_mask = 16'hF0AA;
defparam \halt_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N20
cycloneive_lcell_comb \imemload_id~0 (
// Equation(s):
// imemload_id = (ifid_en1 & (ramiframload_31)) # (!ifid_en1 & ((\prif.imemload_id [31])))

	.dataa(gnd),
	.datab(ramiframload_31),
	.datac(prifimemload_id_31),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id),
	.cout());
// synopsys translate_off
defparam \imemload_id~0 .lut_mask = 16'hCCF0;
defparam \imemload_id~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N22
cycloneive_lcell_comb \imemload_id~1 (
// Equation(s):
// imemload_id1 = (ifid_en1 & (ramiframload_30)) # (!ifid_en1 & ((\prif.imemload_id [30])))

	.dataa(gnd),
	.datab(ramiframload_30),
	.datac(prifimemload_id_30),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id1),
	.cout());
// synopsys translate_off
defparam \imemload_id~1 .lut_mask = 16'hCCF0;
defparam \imemload_id~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N24
cycloneive_lcell_comb \imemload_id~2 (
// Equation(s):
// imemload_id2 = (ifid_en1 & (ramiframload_29)) # (!ifid_en1 & ((\prif.imemload_id [29])))

	.dataa(gnd),
	.datab(ramiframload_29),
	.datac(prifimemload_id_29),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id2),
	.cout());
// synopsys translate_off
defparam \imemload_id~2 .lut_mask = 16'hCCF0;
defparam \imemload_id~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N14
cycloneive_lcell_comb \imemload_id~3 (
// Equation(s):
// imemload_id3 = (ifid_en1 & (ramiframload_27)) # (!ifid_en1 & ((\prif.imemload_id [27])))

	.dataa(gnd),
	.datab(ramiframload_27),
	.datac(prifimemload_id_27),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id3),
	.cout());
// synopsys translate_off
defparam \imemload_id~3 .lut_mask = 16'hCCF0;
defparam \imemload_id~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N16
cycloneive_lcell_comb \imemload_id~4 (
// Equation(s):
// imemload_id4 = (ifid_en1 & (ramiframload_26)) # (!ifid_en1 & ((\prif.imemload_id [26])))

	.dataa(ramiframload_26),
	.datab(gnd),
	.datac(prifimemload_id_26),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id4),
	.cout());
// synopsys translate_off
defparam \imemload_id~4 .lut_mask = 16'hAAF0;
defparam \imemload_id~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N6
cycloneive_lcell_comb \imemload_id~5 (
// Equation(s):
// imemload_id5 = (ifid_en1 & (ramiframload_28)) # (!ifid_en1 & ((\prif.imemload_id [28])))

	.dataa(gnd),
	.datab(ramiframload_28),
	.datac(prifimemload_id_28),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id5),
	.cout());
// synopsys translate_off
defparam \imemload_id~5 .lut_mask = 16'hCCF0;
defparam \imemload_id~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N24
cycloneive_lcell_comb \imemload_id~6 (
// Equation(s):
// imemload_id6 = (ifid_en1 & ((ramiframload_3))) # (!ifid_en1 & (\prif.imemload_id [3]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifimemload_id_3),
	.datad(ramiframload_3),
	.cin(gnd),
	.combout(imemload_id6),
	.cout());
// synopsys translate_off
defparam \imemload_id~6 .lut_mask = 16'hFA50;
defparam \imemload_id~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N8
cycloneive_lcell_comb \imemload_id~7 (
// Equation(s):
// imemload_id7 = (ifid_en1 & (ramiframload_1)) # (!ifid_en1 & ((\prif.imemload_id [1])))

	.dataa(gnd),
	.datab(ramiframload_1),
	.datac(prifimemload_id_1),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id7),
	.cout());
// synopsys translate_off
defparam \imemload_id~7 .lut_mask = 16'hCCF0;
defparam \imemload_id~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N26
cycloneive_lcell_comb \imemload_id~8 (
// Equation(s):
// imemload_id8 = (ifid_en1 & (ramiframload_5)) # (!ifid_en1 & ((\prif.imemload_id [5])))

	.dataa(ifid_en),
	.datab(ramiframload_5),
	.datac(prifimemload_id_5),
	.datad(gnd),
	.cin(gnd),
	.combout(imemload_id8),
	.cout());
// synopsys translate_off
defparam \imemload_id~8 .lut_mask = 16'hD8D8;
defparam \imemload_id~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N28
cycloneive_lcell_comb \imemload_id~9 (
// Equation(s):
// imemload_id9 = (ifid_en1 & ((ramiframload_4))) # (!ifid_en1 & (\prif.imemload_id [4]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifimemload_id_4),
	.datad(ramiframload_4),
	.cin(gnd),
	.combout(imemload_id9),
	.cout());
// synopsys translate_off
defparam \imemload_id~9 .lut_mask = 16'hFA50;
defparam \imemload_id~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N14
cycloneive_lcell_comb \imemload_id~10 (
// Equation(s):
// imemload_id10 = (ifid_en1 & ((ramiframload_2))) # (!ifid_en1 & (\prif.imemload_id [2]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifimemload_id_2),
	.datad(ramiframload_2),
	.cin(gnd),
	.combout(imemload_id10),
	.cout());
// synopsys translate_off
defparam \imemload_id~10 .lut_mask = 16'hFA50;
defparam \imemload_id~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N16
cycloneive_lcell_comb \imemload_id~11 (
// Equation(s):
// imemload_id11 = (ifid_en1 & (ramiframload_0)) # (!ifid_en1 & ((\prif.imemload_id [0])))

	.dataa(ramiframload_0),
	.datab(gnd),
	.datac(prifimemload_id_0),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id11),
	.cout());
// synopsys translate_off
defparam \imemload_id~11 .lut_mask = 16'hAAF0;
defparam \imemload_id~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N30
cycloneive_lcell_comb \imemload_id~12 (
// Equation(s):
// imemload_id12 = (ifid_en1 & (ramiframload_7)) # (!ifid_en1 & ((\prif.imemload_id [7])))

	.dataa(ramiframload_7),
	.datab(gnd),
	.datac(prifimemload_id_7),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id12),
	.cout());
// synopsys translate_off
defparam \imemload_id~12 .lut_mask = 16'hAAF0;
defparam \imemload_id~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N6
cycloneive_lcell_comb \Regwen_ex~0 (
// Equation(s):
// Regwen_ex = (ccifiwait_0 & (((\prif.Regwen_ex~q )))) # (!ccifiwait_0 & ((Selector2) # ((!WideNor0))))

	.dataa(Selector2),
	.datab(ccifiwait_0),
	.datac(prifRegwen_ex),
	.datad(WideNor0),
	.cin(gnd),
	.combout(Regwen_ex),
	.cout());
// synopsys translate_off
defparam \Regwen_ex~0 .lut_mask = 16'hE2F3;
defparam \Regwen_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N24
cycloneive_lcell_comb \rd_ex~0 (
// Equation(s):
// rd_ex = (ccifiwait_0 & (\prif.rd_ex [4])) # (!ccifiwait_0 & ((\prif.imemload_id [15])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrd_ex_4),
	.datad(prifimemload_id_15),
	.cin(gnd),
	.combout(rd_ex),
	.cout());
// synopsys translate_off
defparam \rd_ex~0 .lut_mask = 16'hF5A0;
defparam \rd_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N12
cycloneive_lcell_comb \RegDest_ex~0 (
// Equation(s):
// RegDest_ex = (ccifiwait_0 & (\prif.RegDest_ex [1])) # (!ccifiwait_0 & ((Equal13)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifRegDest_ex_1),
	.datad(Equal13),
	.cin(gnd),
	.combout(RegDest_ex),
	.cout());
// synopsys translate_off
defparam \RegDest_ex~0 .lut_mask = 16'hF3C0;
defparam \RegDest_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N18
cycloneive_lcell_comb \RegDest_ex~1 (
// Equation(s):
// RegDest_ex1 = (ccifiwait_0 & (\prif.RegDest_ex [0])) # (!ccifiwait_0 & ((Selector2)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifRegDest_ex_0),
	.datad(Selector2),
	.cin(gnd),
	.combout(RegDest_ex1),
	.cout());
// synopsys translate_off
defparam \RegDest_ex~1 .lut_mask = 16'hF3C0;
defparam \RegDest_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N18
cycloneive_lcell_comb \rd_ex~1 (
// Equation(s):
// rd_ex1 = (ccifiwait_0 & ((\prif.rd_ex [0]))) # (!ccifiwait_0 & (\prif.imemload_id [11]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_11),
	.datac(prifrd_ex_0),
	.datad(gnd),
	.cin(gnd),
	.combout(rd_ex1),
	.cout());
// synopsys translate_off
defparam \rd_ex~1 .lut_mask = 16'hE4E4;
defparam \rd_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N28
cycloneive_lcell_comb \rd_ex~2 (
// Equation(s):
// rd_ex2 = (ccifiwait_0 & (\prif.rd_ex [1])) # (!ccifiwait_0 & ((\prif.imemload_id [12])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifrd_ex_1),
	.datad(prifimemload_id_12),
	.cin(gnd),
	.combout(rd_ex2),
	.cout());
// synopsys translate_off
defparam \rd_ex~2 .lut_mask = 16'hF3C0;
defparam \rd_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N6
cycloneive_lcell_comb \rd_ex~3 (
// Equation(s):
// rd_ex3 = (ccifiwait_0 & (\prif.rd_ex [2])) # (!ccifiwait_0 & ((\prif.imemload_id [13])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrd_ex_2),
	.datad(prifimemload_id_13),
	.cin(gnd),
	.combout(rd_ex3),
	.cout());
// synopsys translate_off
defparam \rd_ex~3 .lut_mask = 16'hF5A0;
defparam \rd_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N2
cycloneive_lcell_comb \rd_ex~4 (
// Equation(s):
// rd_ex4 = (ccifiwait_0 & (\prif.rd_ex [3])) # (!ccifiwait_0 & ((\prif.imemload_id [14])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifrd_ex_3),
	.datad(prifimemload_id_14),
	.cin(gnd),
	.combout(rd_ex4),
	.cout());
// synopsys translate_off
defparam \rd_ex~4 .lut_mask = 16'hF5A0;
defparam \rd_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N8
cycloneive_lcell_comb \imemload_id~13 (
// Equation(s):
// imemload_id13 = (ifid_en1 & ((ramiframload_17))) # (!ifid_en1 & (\prif.imemload_id [17]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifimemload_id_17),
	.datad(ramiframload_17),
	.cin(gnd),
	.combout(imemload_id13),
	.cout());
// synopsys translate_off
defparam \imemload_id~13 .lut_mask = 16'hFA50;
defparam \imemload_id~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N14
cycloneive_lcell_comb \imemload_id~14 (
// Equation(s):
// imemload_id14 = (ifid_en1 & (ramiframload_16)) # (!ifid_en1 & ((\prif.imemload_id [16])))

	.dataa(gnd),
	.datab(ramiframload_16),
	.datac(prifimemload_id_16),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id14),
	.cout());
// synopsys translate_off
defparam \imemload_id~14 .lut_mask = 16'hCCF0;
defparam \imemload_id~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N8
cycloneive_lcell_comb \imemload_id~15 (
// Equation(s):
// imemload_id15 = (ifid_en1 & (ramiframload_19)) # (!ifid_en1 & ((\prif.imemload_id [19])))

	.dataa(ramiframload_19),
	.datab(gnd),
	.datac(prifimemload_id_19),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id15),
	.cout());
// synopsys translate_off
defparam \imemload_id~15 .lut_mask = 16'hAAF0;
defparam \imemload_id~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N0
cycloneive_lcell_comb \imemload_id~16 (
// Equation(s):
// imemload_id16 = (ifid_en1 & ((ramiframload_18))) # (!ifid_en1 & (\prif.imemload_id [18]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifimemload_id_18),
	.datad(ramiframload_18),
	.cin(gnd),
	.combout(imemload_id16),
	.cout());
// synopsys translate_off
defparam \imemload_id~16 .lut_mask = 16'hFA50;
defparam \imemload_id~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N4
cycloneive_lcell_comb \imemload_id~17 (
// Equation(s):
// imemload_id17 = (ifid_en1 & (ramiframload_20)) # (!ifid_en1 & ((\prif.imemload_id [20])))

	.dataa(ramiframload_20),
	.datab(gnd),
	.datac(prifimemload_id_20),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id17),
	.cout());
// synopsys translate_off
defparam \imemload_id~17 .lut_mask = 16'hAAF0;
defparam \imemload_id~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y31_N0
cycloneive_lcell_comb \dataScr_mem~0 (
// Equation(s):
// dataScr_mem = (exmem_en & ((\prif.dataScr_ex [0]))) # (!exmem_en & (\prif.dataScr_mem [0]))

	.dataa(gnd),
	.datab(exmem_en),
	.datac(prifdataScr_mem_0),
	.datad(prifdataScr_ex_0),
	.cin(gnd),
	.combout(dataScr_mem),
	.cout());
// synopsys translate_off
defparam \dataScr_mem~0 .lut_mask = 16'hFC30;
defparam \dataScr_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N28
cycloneive_lcell_comb \dataScr_mem~1 (
// Equation(s):
// dataScr_mem1 = (exmem_en & ((\prif.dataScr_ex [1]))) # (!exmem_en & (\prif.dataScr_mem [1]))

	.dataa(exmem_en),
	.datab(gnd),
	.datac(prifdataScr_mem_1),
	.datad(prifdataScr_ex_1),
	.cin(gnd),
	.combout(dataScr_mem1),
	.cout());
// synopsys translate_off
defparam \dataScr_mem~1 .lut_mask = 16'hFA50;
defparam \dataScr_mem~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N28
cycloneive_lcell_comb \prif.pc_mem[1]~4 (
// Equation(s):
// prifpc_mem_110 = (\prif.pc_mem[15]~0_combout  & ((\prif.pc_mem [1]))) # (!\prif.pc_mem[15]~0_combout  & (\prif.pc_ex [1]))

	.dataa(prifpc_ex_1),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_1),
	.datad(gnd),
	.cin(gnd),
	.combout(prifpc_mem_110),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[1]~4 .lut_mask = 16'hE2E2;
defparam \prif.pc_mem[1]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N28
cycloneive_lcell_comb \imemload_id~18 (
// Equation(s):
// imemload_id18 = (ifid_en1 & (ramiframload_22)) # (!ifid_en1 & ((\prif.imemload_id [22])))

	.dataa(ramiframload_22),
	.datab(gnd),
	.datac(prifimemload_id_22),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id18),
	.cout());
// synopsys translate_off
defparam \imemload_id~18 .lut_mask = 16'hAAF0;
defparam \imemload_id~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N26
cycloneive_lcell_comb \imemload_id~19 (
// Equation(s):
// imemload_id19 = (ifid_en1 & (ramiframload_21)) # (!ifid_en1 & ((\prif.imemload_id [21])))

	.dataa(ifid_en),
	.datab(ramiframload_21),
	.datac(prifimemload_id_21),
	.datad(gnd),
	.cin(gnd),
	.combout(imemload_id19),
	.cout());
// synopsys translate_off
defparam \imemload_id~19 .lut_mask = 16'hD8D8;
defparam \imemload_id~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N2
cycloneive_lcell_comb \imemload_id~20 (
// Equation(s):
// imemload_id20 = (ifid_en1 & ((ramiframload_24))) # (!ifid_en1 & (\prif.imemload_id [24]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifimemload_id_24),
	.datad(ramiframload_24),
	.cin(gnd),
	.combout(imemload_id20),
	.cout());
// synopsys translate_off
defparam \imemload_id~20 .lut_mask = 16'hFA50;
defparam \imemload_id~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N0
cycloneive_lcell_comb \imemload_id~21 (
// Equation(s):
// imemload_id21 = (ifid_en1 & ((ramiframload_23))) # (!ifid_en1 & (\prif.imemload_id [23]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifimemload_id_23),
	.datad(ramiframload_23),
	.cin(gnd),
	.combout(imemload_id21),
	.cout());
// synopsys translate_off
defparam \imemload_id~21 .lut_mask = 16'hFA50;
defparam \imemload_id~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N12
cycloneive_lcell_comb \imemload_id~22 (
// Equation(s):
// imemload_id22 = (ifid_en1 & (ramiframload_25)) # (!ifid_en1 & ((\prif.imemload_id [25])))

	.dataa(gnd),
	.datab(ramiframload_25),
	.datac(prifimemload_id_25),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id22),
	.cout());
// synopsys translate_off
defparam \imemload_id~22 .lut_mask = 16'hCCF0;
defparam \imemload_id~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N12
cycloneive_lcell_comb \opcode_ex~5 (
// Equation(s):
// opcode_ex5 = (ccifiwait_0 & (\prif.opcode_ex [3])) # (!ccifiwait_0 & ((\prif.imemload_id [29])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifopcode_ex_3),
	.datad(prifimemload_id_29),
	.cin(gnd),
	.combout(opcode_ex5),
	.cout());
// synopsys translate_off
defparam \opcode_ex~5 .lut_mask = 16'hF3C0;
defparam \opcode_ex~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N18
cycloneive_lcell_comb \imemload_id~23 (
// Equation(s):
// imemload_id23 = (ifid_en1 & (ramiframload_6)) # (!ifid_en1 & ((\prif.imemload_id [6])))

	.dataa(ramiframload_6),
	.datab(gnd),
	.datac(prifimemload_id_6),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id23),
	.cout());
// synopsys translate_off
defparam \imemload_id~23 .lut_mask = 16'hAAF0;
defparam \imemload_id~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N26
cycloneive_lcell_comb \prif.pc_mem[0]~5 (
// Equation(s):
// prifpc_mem_01 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [0])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [0])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_0),
	.datad(prifpc_ex_0),
	.cin(gnd),
	.combout(prifpc_mem_01),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[0]~5 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[0]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N8
cycloneive_lcell_comb \prif.pc_mem[3]~6 (
// Equation(s):
// prifpc_mem_32 = (\prif.pc_mem[15]~0_combout  & ((\prif.pc_mem [3]))) # (!\prif.pc_mem[15]~0_combout  & (\prif.pc_ex [3]))

	.dataa(prifpc_ex_3),
	.datab(gnd),
	.datac(prifpc_mem_3),
	.datad(prifpc_mem_151),
	.cin(gnd),
	.combout(prifpc_mem_32),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[3]~6 .lut_mask = 16'hF0AA;
defparam \prif.pc_mem[3]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N4
cycloneive_lcell_comb \imemload_id~24 (
// Equation(s):
// imemload_id24 = (ifid_en1 & (ramiframload_9)) # (!ifid_en1 & ((\prif.imemload_id [9])))

	.dataa(gnd),
	.datab(ramiframload_9),
	.datac(prifimemload_id_9),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id24),
	.cout());
// synopsys translate_off
defparam \imemload_id~24 .lut_mask = 16'hCCF0;
defparam \imemload_id~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N24
cycloneive_lcell_comb \imemload_id~25 (
// Equation(s):
// imemload_id25 = (ifid_en1 & (ramiframload_8)) # (!ifid_en1 & ((\prif.imemload_id [8])))

	.dataa(ifid_en),
	.datab(ramiframload_8),
	.datac(prifimemload_id_8),
	.datad(gnd),
	.cin(gnd),
	.combout(imemload_id25),
	.cout());
// synopsys translate_off
defparam \imemload_id~25 .lut_mask = 16'hD8D8;
defparam \imemload_id~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N26
cycloneive_lcell_comb \prif.pc_mem[2]~7 (
// Equation(s):
// prifpc_mem_210 = (\prif.pc_mem[15]~0_combout  & ((\prif.pc_mem [2]))) # (!\prif.pc_mem[15]~0_combout  & (\prif.pc_ex [2]))

	.dataa(prifpc_ex_2),
	.datab(gnd),
	.datac(prifpc_mem_2),
	.datad(prifpc_mem_151),
	.cin(gnd),
	.combout(prifpc_mem_210),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[2]~7 .lut_mask = 16'hF0AA;
defparam \prif.pc_mem[2]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y27_N24
cycloneive_lcell_comb \prif.pc_mem[4]~8 (
// Equation(s):
// prifpc_mem_41 = (\prif.pc_mem[15]~0_combout  & ((\prif.pc_mem [4]))) # (!\prif.pc_mem[15]~0_combout  & (\prif.pc_ex [4]))

	.dataa(gnd),
	.datab(prifpc_ex_4),
	.datac(prifpc_mem_4),
	.datad(prifpc_mem_151),
	.cin(gnd),
	.combout(prifpc_mem_41),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[4]~8 .lut_mask = 16'hF0CC;
defparam \prif.pc_mem[4]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N2
cycloneive_lcell_comb \imemload_id~26 (
// Equation(s):
// imemload_id26 = (ifid_en1 & ((ramiframload_10))) # (!ifid_en1 & (\prif.imemload_id [10]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifimemload_id_10),
	.datad(ramiframload_10),
	.cin(gnd),
	.combout(imemload_id26),
	.cout());
// synopsys translate_off
defparam \imemload_id~26 .lut_mask = 16'hFA50;
defparam \imemload_id~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N18
cycloneive_lcell_comb \imemload_id~27 (
// Equation(s):
// imemload_id27 = (ifid_en1 & (ramiframload_15)) # (!ifid_en1 & ((\prif.imemload_id [15])))

	.dataa(ramiframload_15),
	.datab(gnd),
	.datac(prifimemload_id_15),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id27),
	.cout());
// synopsys translate_off
defparam \imemload_id~27 .lut_mask = 16'hAAF0;
defparam \imemload_id~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N10
cycloneive_lcell_comb \prif.pc_mem[5]~9 (
// Equation(s):
// prifpc_mem_51 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [5])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [5])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_5),
	.datad(prifpc_ex_5),
	.cin(gnd),
	.combout(prifpc_mem_51),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[5]~9 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[5]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N26
cycloneive_lcell_comb \prif.pc_mem[15]~10 (
// Equation(s):
// prifpc_mem_152 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [15])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [15])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_15),
	.datad(prifpc_ex_15),
	.cin(gnd),
	.combout(prifpc_mem_152),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[15]~10 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[15]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N4
cycloneive_lcell_comb \imemload_id~28 (
// Equation(s):
// imemload_id28 = (ifid_en1 & (ramiframload_14)) # (!ifid_en1 & ((\prif.imemload_id [14])))

	.dataa(ifid_en),
	.datab(ramiframload_14),
	.datac(prifimemload_id_14),
	.datad(gnd),
	.cin(gnd),
	.combout(imemload_id28),
	.cout());
// synopsys translate_off
defparam \imemload_id~28 .lut_mask = 16'hD8D8;
defparam \imemload_id~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N18
cycloneive_lcell_comb \prif.pc_mem[14]~11 (
// Equation(s):
// prifpc_mem_141 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [14])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [14])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_14),
	.datad(prifpc_ex_14),
	.cin(gnd),
	.combout(prifpc_mem_141),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[14]~11 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[14]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N4
cycloneive_lcell_comb \imemload_id~29 (
// Equation(s):
// imemload_id29 = (ifid_en1 & (ramiframload_13)) # (!ifid_en1 & ((\prif.imemload_id [13])))

	.dataa(gnd),
	.datab(ramiframload_13),
	.datac(prifimemload_id_13),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id29),
	.cout());
// synopsys translate_off
defparam \imemload_id~29 .lut_mask = 16'hCCF0;
defparam \imemload_id~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N8
cycloneive_lcell_comb \prif.pc_mem[13]~12 (
// Equation(s):
// prifpc_mem_131 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [13])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [13])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_13),
	.datad(prifpc_ex_13),
	.cin(gnd),
	.combout(prifpc_mem_131),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[13]~12 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[13]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N26
cycloneive_lcell_comb \imemload_id~30 (
// Equation(s):
// imemload_id30 = (ifid_en1 & (ramiframload_12)) # (!ifid_en1 & ((\prif.imemload_id [12])))

	.dataa(gnd),
	.datab(ramiframload_12),
	.datac(prifimemload_id_12),
	.datad(ifid_en),
	.cin(gnd),
	.combout(imemload_id30),
	.cout());
// synopsys translate_off
defparam \imemload_id~30 .lut_mask = 16'hCCF0;
defparam \imemload_id~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N16
cycloneive_lcell_comb \prif.pc_mem[12]~13 (
// Equation(s):
// prifpc_mem_121 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [12])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [12])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_12),
	.datad(prifpc_ex_12),
	.cin(gnd),
	.combout(prifpc_mem_121),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[12]~13 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[12]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N18
cycloneive_lcell_comb \imemload_id~31 (
// Equation(s):
// imemload_id31 = (ifid_en1 & ((ramiframload_11))) # (!ifid_en1 & (\prif.imemload_id [11]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifimemload_id_11),
	.datad(ramiframload_11),
	.cin(gnd),
	.combout(imemload_id31),
	.cout());
// synopsys translate_off
defparam \imemload_id~31 .lut_mask = 16'hFA50;
defparam \imemload_id~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N14
cycloneive_lcell_comb \prif.pc_mem[11]~14 (
// Equation(s):
// prifpc_mem_111 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [11])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [11])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_11),
	.datad(prifpc_ex_11),
	.cin(gnd),
	.combout(prifpc_mem_111),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[11]~14 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[11]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N24
cycloneive_lcell_comb \prif.pc_mem[10]~15 (
// Equation(s):
// prifpc_mem_101 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [10])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [10])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_10),
	.datad(prifpc_ex_10),
	.cin(gnd),
	.combout(prifpc_mem_101),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[10]~15 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[10]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N0
cycloneive_lcell_comb \prif.pc_mem[9]~16 (
// Equation(s):
// prifpc_mem_91 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [9])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [9])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_9),
	.datad(prifpc_ex_9),
	.cin(gnd),
	.combout(prifpc_mem_91),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[9]~16 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[9]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N2
cycloneive_lcell_comb \prif.pc_mem[6]~17 (
// Equation(s):
// prifpc_mem_61 = (\prif.pc_mem[15]~0_combout  & ((\prif.pc_mem [6]))) # (!\prif.pc_mem[15]~0_combout  & (\prif.pc_ex [6]))

	.dataa(prifpc_ex_6),
	.datab(gnd),
	.datac(prifpc_mem_6),
	.datad(prifpc_mem_151),
	.cin(gnd),
	.combout(prifpc_mem_61),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[6]~17 .lut_mask = 16'hF0AA;
defparam \prif.pc_mem[6]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N20
cycloneive_lcell_comb \prif.pc_mem[27]~18 (
// Equation(s):
// prifpc_mem_271 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [27])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [27])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_27),
	.datad(prifpc_ex_27),
	.cin(gnd),
	.combout(prifpc_mem_271),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[27]~18 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[27]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N18
cycloneive_lcell_comb \prif.pc_mem[23]~19 (
// Equation(s):
// prifpc_mem_231 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [23])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [23])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_23),
	.datad(prifpc_ex_23),
	.cin(gnd),
	.combout(prifpc_mem_231),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[23]~19 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[23]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N16
cycloneive_lcell_comb \prif.pc_mem[18]~20 (
// Equation(s):
// prifpc_mem_181 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [18])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [18])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_18),
	.datad(prifpc_ex_18),
	.cin(gnd),
	.combout(prifpc_mem_181),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[18]~20 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[18]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N30
cycloneive_lcell_comb \prif.pc_mem[24]~21 (
// Equation(s):
// prifpc_mem_241 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [24])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [24])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_24),
	.datad(prifpc_ex_24),
	.cin(gnd),
	.combout(prifpc_mem_241),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[24]~21 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[24]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N20
cycloneive_lcell_comb \prif.pc_mem[16]~22 (
// Equation(s):
// prifpc_mem_161 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [16])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [16])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_16),
	.datad(prifpc_ex_16),
	.cin(gnd),
	.combout(prifpc_mem_161),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[16]~22 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[16]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N8
cycloneive_lcell_comb \prif.pc_mem[19]~23 (
// Equation(s):
// prifpc_mem_191 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [19])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [19])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_19),
	.datad(prifpc_ex_19),
	.cin(gnd),
	.combout(prifpc_mem_191),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[19]~23 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[19]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N22
cycloneive_lcell_comb \prif.pc_mem[17]~24 (
// Equation(s):
// prifpc_mem_171 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [17])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [17])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_17),
	.datad(prifpc_ex_17),
	.cin(gnd),
	.combout(prifpc_mem_171),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[17]~24 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[17]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N4
cycloneive_lcell_comb \prif.pc_mem[21]~25 (
// Equation(s):
// prifpc_mem_211 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [21])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [21])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_21),
	.datad(prifpc_ex_21),
	.cin(gnd),
	.combout(prifpc_mem_211),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[21]~25 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[21]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N14
cycloneive_lcell_comb \prif.pc_mem[20]~26 (
// Equation(s):
// prifpc_mem_201 = (\prif.pc_mem[15]~0_combout  & ((\prif.pc_mem [20]))) # (!\prif.pc_mem[15]~0_combout  & (\prif.pc_ex [20]))

	.dataa(gnd),
	.datab(prifpc_ex_20),
	.datac(prifpc_mem_20),
	.datad(prifpc_mem_151),
	.cin(gnd),
	.combout(prifpc_mem_201),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[20]~26 .lut_mask = 16'hF0CC;
defparam \prif.pc_mem[20]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N6
cycloneive_lcell_comb \prif.pc_mem[26]~27 (
// Equation(s):
// prifpc_mem_261 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [26])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [26])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_26),
	.datad(prifpc_ex_26),
	.cin(gnd),
	.combout(prifpc_mem_261),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[26]~27 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[26]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N20
cycloneive_lcell_comb \prif.pc_mem[8]~28 (
// Equation(s):
// prifpc_mem_81 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [8])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [8])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_8),
	.datad(prifpc_ex_8),
	.cin(gnd),
	.combout(prifpc_mem_81),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[8]~28 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[8]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N6
cycloneive_lcell_comb \prif.pc_mem[7]~29 (
// Equation(s):
// prifpc_mem_71 = (\prif.pc_mem[15]~0_combout  & ((\prif.pc_mem [7]))) # (!\prif.pc_mem[15]~0_combout  & (\prif.pc_ex [7]))

	.dataa(prifpc_ex_7),
	.datab(gnd),
	.datac(prifpc_mem_7),
	.datad(prifpc_mem_151),
	.cin(gnd),
	.combout(prifpc_mem_71),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[7]~29 .lut_mask = 16'hF0AA;
defparam \prif.pc_mem[7]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N22
cycloneive_lcell_comb \prif.pc_mem[22]~30 (
// Equation(s):
// prifpc_mem_221 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [22])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [22])))

	.dataa(prifpc_mem_151),
	.datab(gnd),
	.datac(prifpc_mem_22),
	.datad(prifpc_ex_22),
	.cin(gnd),
	.combout(prifpc_mem_221),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[22]~30 .lut_mask = 16'hF5A0;
defparam \prif.pc_mem[22]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N2
cycloneive_lcell_comb \prif.pc_mem[25]~31 (
// Equation(s):
// prifpc_mem_251 = (\prif.pc_mem[15]~0_combout  & (\prif.pc_mem [25])) # (!\prif.pc_mem[15]~0_combout  & ((\prif.pc_ex [25])))

	.dataa(gnd),
	.datab(prifpc_mem_151),
	.datac(prifpc_mem_25),
	.datad(prifpc_ex_25),
	.cin(gnd),
	.combout(prifpc_mem_251),
	.cout());
// synopsys translate_off
defparam \prif.pc_mem[25]~31 .lut_mask = 16'hF3C0;
defparam \prif.pc_mem[25]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N30
cycloneive_lcell_comb \instr_ex~1 (
// Equation(s):
// instr_ex1 = (ccifiwait_0 & (\prif.instr_ex [3])) # (!ccifiwait_0 & ((\prif.imemload_id [3])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_3),
	.datad(prifimemload_id_3),
	.cin(gnd),
	.combout(instr_ex1),
	.cout());
// synopsys translate_off
defparam \instr_ex~1 .lut_mask = 16'hF5A0;
defparam \instr_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N10
cycloneive_lcell_comb \instr_ex~2 (
// Equation(s):
// instr_ex2 = (ccifiwait_0 & (\prif.instr_ex [5])) # (!ccifiwait_0 & ((\prif.imemload_id [5])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifinstr_ex_5),
	.datad(prifimemload_id_5),
	.cin(gnd),
	.combout(instr_ex2),
	.cout());
// synopsys translate_off
defparam \instr_ex~2 .lut_mask = 16'hF3C0;
defparam \instr_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N28
cycloneive_lcell_comb \instr_ex~3 (
// Equation(s):
// instr_ex3 = (ccifiwait_0 & (\prif.instr_ex [4])) # (!ccifiwait_0 & ((\prif.imemload_id [4])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifinstr_ex_4),
	.datad(prifimemload_id_4),
	.cin(gnd),
	.combout(instr_ex3),
	.cout());
// synopsys translate_off
defparam \instr_ex~3 .lut_mask = 16'hF3C0;
defparam \instr_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N6
cycloneive_lcell_comb \instr_ex~4 (
// Equation(s):
// instr_ex4 = (ccifiwait_0 & (\prif.instr_ex [2])) # (!ccifiwait_0 & ((\prif.imemload_id [2])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifinstr_ex_2),
	.datad(prifimemload_id_2),
	.cin(gnd),
	.combout(instr_ex4),
	.cout());
// synopsys translate_off
defparam \instr_ex~4 .lut_mask = 16'hF3C0;
defparam \instr_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N0
cycloneive_lcell_comb \instr_ex~5 (
// Equation(s):
// instr_ex5 = (ccifiwait_0 & (\prif.instr_ex [1])) # (!ccifiwait_0 & ((\prif.imemload_id [1])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_1),
	.datad(prifimemload_id_1),
	.cin(gnd),
	.combout(instr_ex5),
	.cout());
// synopsys translate_off
defparam \instr_ex~5 .lut_mask = 16'hF5A0;
defparam \instr_ex~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y28_N2
cycloneive_lcell_comb \instr_ex~6 (
// Equation(s):
// instr_ex6 = (ccifiwait_0 & (\prif.instr_ex [0])) # (!ccifiwait_0 & ((\prif.imemload_id [0])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_0),
	.datad(prifimemload_id_0),
	.cin(gnd),
	.combout(instr_ex6),
	.cout());
// synopsys translate_off
defparam \instr_ex~6 .lut_mask = 16'hF5A0;
defparam \instr_ex~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N28
cycloneive_lcell_comb \PCScr_ex~3 (
// Equation(s):
// PCScr_ex = (ccifiwait_0 & (((\prif.PCScr_ex [0])))) # (!ccifiwait_0 & (((!ALUScr_ex2)) # (!\PCScr_ex~2_combout )))

	.dataa(ccifiwait_0),
	.datab(\PCScr_ex~2_combout ),
	.datac(prifPCScr_ex_0),
	.datad(ALUScr_ex2),
	.cin(gnd),
	.combout(PCScr_ex),
	.cout());
// synopsys translate_off
defparam \PCScr_ex~3 .lut_mask = 16'hB1F5;
defparam \PCScr_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N30
cycloneive_lcell_comb \pc_ex~0 (
// Equation(s):
// pc_ex = (ccifiwait_0 & (\prif.pc_ex [1])) # (!ccifiwait_0 & ((\prif.pc_id [1])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifpc_ex_1),
	.datad(prifpc_id_1),
	.cin(gnd),
	.combout(pc_ex),
	.cout());
// synopsys translate_off
defparam \pc_ex~0 .lut_mask = 16'hF3C0;
defparam \pc_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N4
cycloneive_lcell_comb \PCScr_ex~4 (
// Equation(s):
// PCScr_ex1 = (ccifiwait_0 & (\prif.PCScr_ex [1])) # (!ccifiwait_0 & ((\PCScr_ex~5_combout )))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifPCScr_ex_1),
	.datad(\PCScr_ex~5_combout ),
	.cin(gnd),
	.combout(PCScr_ex1),
	.cout());
// synopsys translate_off
defparam \PCScr_ex~4 .lut_mask = 16'hF5A0;
defparam \PCScr_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N16
cycloneive_lcell_comb \pc_ex~1 (
// Equation(s):
// pc_ex1 = (ccifiwait_0 & ((\prif.pc_ex [0]))) # (!ccifiwait_0 & (\prif.pc_id [0]))

	.dataa(prifpc_id_0),
	.datab(ccifiwait_0),
	.datac(prifpc_ex_0),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_ex1),
	.cout());
// synopsys translate_off
defparam \pc_ex~1 .lut_mask = 16'hE2E2;
defparam \pc_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N20
cycloneive_lcell_comb \pc_ex~2 (
// Equation(s):
// pc_ex2 = (ccifiwait_0 & (\prif.pc_ex [3])) # (!ccifiwait_0 & ((\prif.pc_id [3])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifpc_ex_3),
	.datad(prifpc_id_3),
	.cin(gnd),
	.combout(pc_ex2),
	.cout());
// synopsys translate_off
defparam \pc_ex~2 .lut_mask = 16'hF3C0;
defparam \pc_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N8
cycloneive_lcell_comb \pc_ex~3 (
// Equation(s):
// pc_ex3 = (ccifiwait_0 & (\prif.pc_ex [2])) # (!ccifiwait_0 & ((\prif.pc_id [2])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_2),
	.datad(prifpc_id_2),
	.cin(gnd),
	.combout(pc_ex3),
	.cout());
// synopsys translate_off
defparam \pc_ex~3 .lut_mask = 16'hF5A0;
defparam \pc_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N0
cycloneive_lcell_comb \pc_ex~4 (
// Equation(s):
// pc_ex4 = (ccifiwait_0 & ((\prif.pc_ex [5]))) # (!ccifiwait_0 & (\prif.pc_id [5]))

	.dataa(ccifiwait_0),
	.datab(prifpc_id_5),
	.datac(prifpc_ex_5),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_ex4),
	.cout());
// synopsys translate_off
defparam \pc_ex~4 .lut_mask = 16'hE4E4;
defparam \pc_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N22
cycloneive_lcell_comb \pc_ex~5 (
// Equation(s):
// pc_ex5 = (ccifiwait_0 & (\prif.pc_ex [4])) # (!ccifiwait_0 & ((\prif.pc_id [4])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_4),
	.datad(prifpc_id_4),
	.cin(gnd),
	.combout(pc_ex5),
	.cout());
// synopsys translate_off
defparam \pc_ex~5 .lut_mask = 16'hF5A0;
defparam \pc_ex~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N30
cycloneive_lcell_comb \pc_ex~6 (
// Equation(s):
// pc_ex6 = (ccifiwait_0 & (\prif.pc_ex [7])) # (!ccifiwait_0 & ((\prif.pc_id [7])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_7),
	.datad(prifpc_id_7),
	.cin(gnd),
	.combout(pc_ex6),
	.cout());
// synopsys translate_off
defparam \pc_ex~6 .lut_mask = 16'hF5A0;
defparam \pc_ex~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N12
cycloneive_lcell_comb \pc_ex~7 (
// Equation(s):
// pc_ex7 = (ccifiwait_0 & (\prif.pc_ex [6])) # (!ccifiwait_0 & ((\prif.pc_id [6])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_6),
	.datad(prifpc_id_6),
	.cin(gnd),
	.combout(pc_ex7),
	.cout());
// synopsys translate_off
defparam \pc_ex~7 .lut_mask = 16'hF5A0;
defparam \pc_ex~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N10
cycloneive_lcell_comb \pc_ex~8 (
// Equation(s):
// pc_ex8 = (ccifiwait_0 & (\prif.pc_ex [9])) # (!ccifiwait_0 & ((\prif.pc_id [9])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_9),
	.datad(prifpc_id_9),
	.cin(gnd),
	.combout(pc_ex8),
	.cout());
// synopsys translate_off
defparam \pc_ex~8 .lut_mask = 16'hF5A0;
defparam \pc_ex~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y33_N16
cycloneive_lcell_comb \pc_ex~9 (
// Equation(s):
// pc_ex9 = (ccifiwait_0 & ((\prif.pc_ex [8]))) # (!ccifiwait_0 & (\prif.pc_id [8]))

	.dataa(ccifiwait_0),
	.datab(prifpc_id_8),
	.datac(prifpc_ex_8),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_ex9),
	.cout());
// synopsys translate_off
defparam \pc_ex~9 .lut_mask = 16'hE4E4;
defparam \pc_ex~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y23_N6
cycloneive_lcell_comb \instr_ex~7 (
// Equation(s):
// instr_ex7 = (ccifiwait_0 & ((\prif.instr_ex [7]))) # (!ccifiwait_0 & (\prif.imemload_id [7]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_7),
	.datac(prifinstr_ex_7),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_ex7),
	.cout());
// synopsys translate_off
defparam \instr_ex~7 .lut_mask = 16'hE4E4;
defparam \instr_ex~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N6
cycloneive_lcell_comb \instr_ex~8 (
// Equation(s):
// instr_ex8 = (ccifiwait_0 & (\prif.instr_ex [6])) # (!ccifiwait_0 & ((\prif.imemload_id [6])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_6),
	.datad(prifimemload_id_6),
	.cin(gnd),
	.combout(instr_ex8),
	.cout());
// synopsys translate_off
defparam \instr_ex~8 .lut_mask = 16'hF5A0;
defparam \instr_ex~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N28
cycloneive_lcell_comb \pc_ex~10 (
// Equation(s):
// pc_ex10 = (ccifiwait_0 & (\prif.pc_ex [11])) # (!ccifiwait_0 & ((\prif.pc_id [11])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_11),
	.datad(prifpc_id_11),
	.cin(gnd),
	.combout(pc_ex10),
	.cout());
// synopsys translate_off
defparam \pc_ex~10 .lut_mask = 16'hF5A0;
defparam \pc_ex~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N2
cycloneive_lcell_comb \pc_ex~11 (
// Equation(s):
// pc_ex11 = (ccifiwait_0 & (\prif.pc_ex [10])) # (!ccifiwait_0 & ((\prif.pc_id [10])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_10),
	.datad(prifpc_id_10),
	.cin(gnd),
	.combout(pc_ex11),
	.cout());
// synopsys translate_off
defparam \pc_ex~11 .lut_mask = 16'hF5A0;
defparam \pc_ex~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N8
cycloneive_lcell_comb \instr_ex~9 (
// Equation(s):
// instr_ex9 = (ccifiwait_0 & (\prif.instr_ex [9])) # (!ccifiwait_0 & ((\prif.imemload_id [9])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifinstr_ex_9),
	.datad(prifimemload_id_9),
	.cin(gnd),
	.combout(instr_ex9),
	.cout());
// synopsys translate_off
defparam \instr_ex~9 .lut_mask = 16'hF3C0;
defparam \instr_ex~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N12
cycloneive_lcell_comb \instr_ex~10 (
// Equation(s):
// instr_ex10 = (ccifiwait_0 & (\prif.instr_ex [8])) # (!ccifiwait_0 & ((\prif.imemload_id [8])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_8),
	.datad(prifimemload_id_8),
	.cin(gnd),
	.combout(instr_ex10),
	.cout());
// synopsys translate_off
defparam \instr_ex~10 .lut_mask = 16'hF5A0;
defparam \instr_ex~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N0
cycloneive_lcell_comb \pc_ex~12 (
// Equation(s):
// pc_ex12 = (ccifiwait_0 & (\prif.pc_ex [13])) # (!ccifiwait_0 & ((\prif.pc_id [13])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_13),
	.datad(prifpc_id_13),
	.cin(gnd),
	.combout(pc_ex12),
	.cout());
// synopsys translate_off
defparam \pc_ex~12 .lut_mask = 16'hF5A0;
defparam \pc_ex~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N18
cycloneive_lcell_comb \pc_ex~13 (
// Equation(s):
// pc_ex13 = (ccifiwait_0 & (\prif.pc_ex [12])) # (!ccifiwait_0 & ((\prif.pc_id [12])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_12),
	.datad(prifpc_id_12),
	.cin(gnd),
	.combout(pc_ex13),
	.cout());
// synopsys translate_off
defparam \pc_ex~13 .lut_mask = 16'hF5A0;
defparam \pc_ex~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N24
cycloneive_lcell_comb \instr_ex~11 (
// Equation(s):
// instr_ex11 = (ccifiwait_0 & ((\prif.instr_ex [11]))) # (!ccifiwait_0 & (\prif.imemload_id [11]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_11),
	.datac(prifinstr_ex_11),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_ex11),
	.cout());
// synopsys translate_off
defparam \instr_ex~11 .lut_mask = 16'hE4E4;
defparam \instr_ex~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N14
cycloneive_lcell_comb \instr_ex~12 (
// Equation(s):
// instr_ex12 = (ccifiwait_0 & (\prif.instr_ex [10])) # (!ccifiwait_0 & ((\prif.imemload_id [10])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifinstr_ex_10),
	.datad(prifimemload_id_10),
	.cin(gnd),
	.combout(instr_ex12),
	.cout());
// synopsys translate_off
defparam \instr_ex~12 .lut_mask = 16'hF3C0;
defparam \instr_ex~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N20
cycloneive_lcell_comb \pc_ex~14 (
// Equation(s):
// pc_ex14 = (ccifiwait_0 & (\prif.pc_ex [15])) # (!ccifiwait_0 & ((\prif.pc_id [15])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_15),
	.datad(prifpc_id_15),
	.cin(gnd),
	.combout(pc_ex14),
	.cout());
// synopsys translate_off
defparam \pc_ex~14 .lut_mask = 16'hF5A0;
defparam \pc_ex~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N30
cycloneive_lcell_comb \pc_ex~15 (
// Equation(s):
// pc_ex15 = (ccifiwait_0 & (\prif.pc_ex [14])) # (!ccifiwait_0 & ((\prif.pc_id [14])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifpc_ex_14),
	.datad(prifpc_id_14),
	.cin(gnd),
	.combout(pc_ex15),
	.cout());
// synopsys translate_off
defparam \pc_ex~15 .lut_mask = 16'hF3C0;
defparam \pc_ex~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N10
cycloneive_lcell_comb \instr_ex~13 (
// Equation(s):
// instr_ex13 = (ccifiwait_0 & (\prif.instr_ex [13])) # (!ccifiwait_0 & ((\prif.imemload_id [13])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_13),
	.datad(prifimemload_id_13),
	.cin(gnd),
	.combout(instr_ex13),
	.cout());
// synopsys translate_off
defparam \instr_ex~13 .lut_mask = 16'hF5A0;
defparam \instr_ex~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N14
cycloneive_lcell_comb \instr_ex~14 (
// Equation(s):
// instr_ex14 = (ccifiwait_0 & (\prif.instr_ex [12])) # (!ccifiwait_0 & ((\prif.imemload_id [12])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifinstr_ex_12),
	.datad(prifimemload_id_12),
	.cin(gnd),
	.combout(instr_ex14),
	.cout());
// synopsys translate_off
defparam \instr_ex~14 .lut_mask = 16'hF3C0;
defparam \instr_ex~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N10
cycloneive_lcell_comb \pc_ex~16 (
// Equation(s):
// pc_ex16 = (ccifiwait_0 & (\prif.pc_ex [23])) # (!ccifiwait_0 & ((\prif.pc_id [23])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_23),
	.datad(prifpc_id_23),
	.cin(gnd),
	.combout(pc_ex16),
	.cout());
// synopsys translate_off
defparam \pc_ex~16 .lut_mask = 16'hF5A0;
defparam \pc_ex~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N8
cycloneive_lcell_comb \pc_ex~17 (
// Equation(s):
// pc_ex17 = (ccifiwait_0 & ((\prif.pc_ex [22]))) # (!ccifiwait_0 & (\prif.pc_id [22]))

	.dataa(prifpc_id_22),
	.datab(ccifiwait_0),
	.datac(prifpc_ex_22),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_ex17),
	.cout());
// synopsys translate_off
defparam \pc_ex~17 .lut_mask = 16'hE2E2;
defparam \pc_ex~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N0
cycloneive_lcell_comb \pc_ex~18 (
// Equation(s):
// pc_ex18 = (ccifiwait_0 & (\prif.pc_ex [21])) # (!ccifiwait_0 & ((\prif.pc_id [21])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_21),
	.datad(prifpc_id_21),
	.cin(gnd),
	.combout(pc_ex18),
	.cout());
// synopsys translate_off
defparam \pc_ex~18 .lut_mask = 16'hF5A0;
defparam \pc_ex~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y31_N0
cycloneive_lcell_comb \pc_ex~19 (
// Equation(s):
// pc_ex19 = (ccifiwait_0 & (\prif.pc_ex [20])) # (!ccifiwait_0 & ((\prif.pc_id [20])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifpc_ex_20),
	.datad(prifpc_id_20),
	.cin(gnd),
	.combout(pc_ex19),
	.cout());
// synopsys translate_off
defparam \pc_ex~19 .lut_mask = 16'hF3C0;
defparam \pc_ex~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N2
cycloneive_lcell_comb \pc_ex~20 (
// Equation(s):
// pc_ex20 = (ccifiwait_0 & (\prif.pc_ex [19])) # (!ccifiwait_0 & ((\prif.pc_id [19])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_19),
	.datad(prifpc_id_19),
	.cin(gnd),
	.combout(pc_ex20),
	.cout());
// synopsys translate_off
defparam \pc_ex~20 .lut_mask = 16'hF5A0;
defparam \pc_ex~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N12
cycloneive_lcell_comb \pc_ex~21 (
// Equation(s):
// pc_ex21 = (ccifiwait_0 & ((\prif.pc_ex [18]))) # (!ccifiwait_0 & (\prif.pc_id [18]))

	.dataa(ccifiwait_0),
	.datab(prifpc_id_18),
	.datac(prifpc_ex_18),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_ex21),
	.cout());
// synopsys translate_off
defparam \pc_ex~21 .lut_mask = 16'hE4E4;
defparam \pc_ex~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N26
cycloneive_lcell_comb \pc_ex~22 (
// Equation(s):
// pc_ex22 = (ccifiwait_0 & (\prif.pc_ex [17])) # (!ccifiwait_0 & ((\prif.pc_id [17])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_17),
	.datad(prifpc_id_17),
	.cin(gnd),
	.combout(pc_ex22),
	.cout());
// synopsys translate_off
defparam \pc_ex~22 .lut_mask = 16'hF5A0;
defparam \pc_ex~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N8
cycloneive_lcell_comb \pc_ex~23 (
// Equation(s):
// pc_ex23 = (ccifiwait_0 & (\prif.pc_ex [16])) # (!ccifiwait_0 & ((\prif.pc_id [16])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_16),
	.datad(prifpc_id_16),
	.cin(gnd),
	.combout(pc_ex23),
	.cout());
// synopsys translate_off
defparam \pc_ex~23 .lut_mask = 16'hF5A0;
defparam \pc_ex~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y31_N30
cycloneive_lcell_comb \instr_ex~15 (
// Equation(s):
// instr_ex15 = (ccifiwait_0 & (\prif.instr_ex [21])) # (!ccifiwait_0 & ((\prif.imemload_id [21])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_21),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(instr_ex15),
	.cout());
// synopsys translate_off
defparam \instr_ex~15 .lut_mask = 16'hF5A0;
defparam \instr_ex~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N20
cycloneive_lcell_comb \instr_ex~16 (
// Equation(s):
// instr_ex16 = (ccifiwait_0 & (\prif.instr_ex [20])) # (!ccifiwait_0 & ((\prif.imemload_id [20])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifinstr_ex_20),
	.datad(prifimemload_id_20),
	.cin(gnd),
	.combout(instr_ex16),
	.cout());
// synopsys translate_off
defparam \instr_ex~16 .lut_mask = 16'hF3C0;
defparam \instr_ex~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N16
cycloneive_lcell_comb \instr_ex~17 (
// Equation(s):
// instr_ex17 = (ccifiwait_0 & (\prif.instr_ex [19])) # (!ccifiwait_0 & ((\prif.imemload_id [19])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_19),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(instr_ex17),
	.cout());
// synopsys translate_off
defparam \instr_ex~17 .lut_mask = 16'hF5A0;
defparam \instr_ex~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N14
cycloneive_lcell_comb \pc_ex~24 (
// Equation(s):
// pc_ex24 = (ccifiwait_0 & (\prif.pc_ex [29])) # (!ccifiwait_0 & ((\prif.pc_id [29])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_29),
	.datad(prifpc_id_29),
	.cin(gnd),
	.combout(pc_ex24),
	.cout());
// synopsys translate_off
defparam \pc_ex~24 .lut_mask = 16'hF5A0;
defparam \pc_ex~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N2
cycloneive_lcell_comb \pc_ex~25 (
// Equation(s):
// pc_ex25 = (ccifiwait_0 & (\prif.pc_ex [28])) # (!ccifiwait_0 & ((\prif.pc_id [28])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifpc_ex_28),
	.datad(prifpc_id_28),
	.cin(gnd),
	.combout(pc_ex25),
	.cout());
// synopsys translate_off
defparam \pc_ex~25 .lut_mask = 16'hF3C0;
defparam \pc_ex~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N10
cycloneive_lcell_comb \pc_ex~26 (
// Equation(s):
// pc_ex26 = (ccifiwait_0 & (\prif.pc_ex [27])) # (!ccifiwait_0 & ((\prif.pc_id [27])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_27),
	.datad(prifpc_id_27),
	.cin(gnd),
	.combout(pc_ex26),
	.cout());
// synopsys translate_off
defparam \pc_ex~26 .lut_mask = 16'hF5A0;
defparam \pc_ex~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y32_N24
cycloneive_lcell_comb \pc_ex~27 (
// Equation(s):
// pc_ex27 = (ccifiwait_0 & (\prif.pc_ex [26])) # (!ccifiwait_0 & ((\prif.pc_id [26])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_26),
	.datad(prifpc_id_26),
	.cin(gnd),
	.combout(pc_ex27),
	.cout());
// synopsys translate_off
defparam \pc_ex~27 .lut_mask = 16'hF5A0;
defparam \pc_ex~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N12
cycloneive_lcell_comb \pc_ex~28 (
// Equation(s):
// pc_ex28 = (ccifiwait_0 & ((\prif.pc_ex [25]))) # (!ccifiwait_0 & (\prif.pc_id [25]))

	.dataa(ccifiwait_0),
	.datab(prifpc_id_25),
	.datac(prifpc_ex_25),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_ex28),
	.cout());
// synopsys translate_off
defparam \pc_ex~28 .lut_mask = 16'hE4E4;
defparam \pc_ex~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N4
cycloneive_lcell_comb \pc_ex~29 (
// Equation(s):
// pc_ex29 = (ccifiwait_0 & (\prif.pc_ex [24])) # (!ccifiwait_0 & ((\prif.pc_id [24])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifpc_ex_24),
	.datad(prifpc_id_24),
	.cin(gnd),
	.combout(pc_ex29),
	.cout());
// synopsys translate_off
defparam \pc_ex~29 .lut_mask = 16'hF5A0;
defparam \pc_ex~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N0
cycloneive_lcell_comb \pc_ex~30 (
// Equation(s):
// pc_ex30 = (ccifiwait_0 & (\prif.pc_ex [31])) # (!ccifiwait_0 & ((\prif.pc_id [31])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifpc_ex_31),
	.datad(prifpc_id_31),
	.cin(gnd),
	.combout(pc_ex30),
	.cout());
// synopsys translate_off
defparam \pc_ex~30 .lut_mask = 16'hF3C0;
defparam \pc_ex~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y34_N14
cycloneive_lcell_comb \pc_ex~31 (
// Equation(s):
// pc_ex31 = (ccifiwait_0 & (\prif.pc_ex [30])) # (!ccifiwait_0 & ((\prif.pc_id [30])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifpc_ex_30),
	.datad(prifpc_id_30),
	.cin(gnd),
	.combout(pc_ex31),
	.cout());
// synopsys translate_off
defparam \pc_ex~31 .lut_mask = 16'hF3C0;
defparam \pc_ex~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N30
cycloneive_lcell_comb \instr_ex~18 (
// Equation(s):
// instr_ex18 = (ccifiwait_0 & ((\prif.instr_ex [18]))) # (!ccifiwait_0 & (\prif.imemload_id [18]))

	.dataa(prifimemload_id_18),
	.datab(gnd),
	.datac(prifinstr_ex_18),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(instr_ex18),
	.cout());
// synopsys translate_off
defparam \instr_ex~18 .lut_mask = 16'hF0AA;
defparam \instr_ex~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N30
cycloneive_lcell_comb \instr_ex~19 (
// Equation(s):
// instr_ex19 = (ccifiwait_0 & (\prif.instr_ex [14])) # (!ccifiwait_0 & ((\prif.imemload_id [14])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_14),
	.datad(prifimemload_id_14),
	.cin(gnd),
	.combout(instr_ex19),
	.cout());
// synopsys translate_off
defparam \instr_ex~19 .lut_mask = 16'hF5A0;
defparam \instr_ex~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N30
cycloneive_lcell_comb \instr_ex~20 (
// Equation(s):
// instr_ex20 = (ccifiwait_0 & (\prif.instr_ex [17])) # (!ccifiwait_0 & ((\prif.imemload_id [17])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_17),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(instr_ex20),
	.cout());
// synopsys translate_off
defparam \instr_ex~20 .lut_mask = 16'hF5A0;
defparam \instr_ex~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N16
cycloneive_lcell_comb \instr_ex~21 (
// Equation(s):
// instr_ex21 = (ccifiwait_0 & ((\prif.instr_ex [16]))) # (!ccifiwait_0 & (\prif.imemload_id [16]))

	.dataa(prifimemload_id_16),
	.datab(gnd),
	.datac(prifinstr_ex_16),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(instr_ex21),
	.cout());
// synopsys translate_off
defparam \instr_ex~21 .lut_mask = 16'hF0AA;
defparam \instr_ex~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N2
cycloneive_lcell_comb \instr_ex~22 (
// Equation(s):
// instr_ex22 = (ccifiwait_0 & ((\prif.instr_ex [23]))) # (!ccifiwait_0 & (\prif.imemload_id [23]))

	.dataa(gnd),
	.datab(prifimemload_id_23),
	.datac(prifinstr_ex_23),
	.datad(ccifiwait_0),
	.cin(gnd),
	.combout(instr_ex22),
	.cout());
// synopsys translate_off
defparam \instr_ex~22 .lut_mask = 16'hF0CC;
defparam \instr_ex~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N24
cycloneive_lcell_comb \instr_ex~23 (
// Equation(s):
// instr_ex23 = (ccifiwait_0 & (\prif.instr_ex [22])) # (!ccifiwait_0 & ((\prif.imemload_id [22])))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifinstr_ex_22),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(instr_ex23),
	.cout());
// synopsys translate_off
defparam \instr_ex~23 .lut_mask = 16'hF3C0;
defparam \instr_ex~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y32_N8
cycloneive_lcell_comb \instr_ex~24 (
// Equation(s):
// instr_ex24 = (ccifiwait_0 & (\prif.instr_ex [25])) # (!ccifiwait_0 & ((\prif.imemload_id [25])))

	.dataa(ccifiwait_0),
	.datab(gnd),
	.datac(prifinstr_ex_25),
	.datad(prifimemload_id_25),
	.cin(gnd),
	.combout(instr_ex24),
	.cout());
// synopsys translate_off
defparam \instr_ex~24 .lut_mask = 16'hF5A0;
defparam \instr_ex~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y33_N28
cycloneive_lcell_comb \instr_ex~25 (
// Equation(s):
// instr_ex25 = (ccifiwait_0 & ((\prif.instr_ex [24]))) # (!ccifiwait_0 & (\prif.imemload_id [24]))

	.dataa(ccifiwait_0),
	.datab(prifimemload_id_24),
	.datac(prifinstr_ex_24),
	.datad(gnd),
	.cin(gnd),
	.combout(instr_ex25),
	.cout());
// synopsys translate_off
defparam \instr_ex~25 .lut_mask = 16'hE4E4;
defparam \instr_ex~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y29_N2
cycloneive_lcell_comb \halt_wb~0 (
// Equation(s):
// halt_wb = (always1 & ((\prif.halt_mem~q ))) # (!always1 & (\prif.halt_wb~q ))

	.dataa(gnd),
	.datab(always1),
	.datac(prifhalt_wb),
	.datad(prifhalt_mem),
	.cin(gnd),
	.combout(halt_wb),
	.cout());
// synopsys translate_off
defparam \halt_wb~0 .lut_mask = 16'hFC30;
defparam \halt_wb~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N20
cycloneive_lcell_comb \dataScr_ex~3 (
// Equation(s):
// dataScr_ex1 = (ccifiwait_0 & (\prif.dataScr_ex [1])) # (!ccifiwait_0 & ((!dataScr_ex)))

	.dataa(gnd),
	.datab(ccifiwait_0),
	.datac(prifdataScr_ex_1),
	.datad(dataScr_ex),
	.cin(gnd),
	.combout(dataScr_ex1),
	.cout());
// synopsys translate_off
defparam \dataScr_ex~3 .lut_mask = 16'hC0F3;
defparam \dataScr_ex~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N8
cycloneive_lcell_comb \pc_id~0 (
// Equation(s):
// pc_id = (ifid_en1 & (pc_1)) # (!ifid_en1 & ((\prif.pc_id [1])))

	.dataa(ifid_en),
	.datab(pc_1),
	.datac(prifpc_id_1),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_id),
	.cout());
// synopsys translate_off
defparam \pc_id~0 .lut_mask = 16'hD8D8;
defparam \pc_id~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N6
cycloneive_lcell_comb \pc_id~1 (
// Equation(s):
// pc_id1 = (ifid_en1 & (pc_0)) # (!ifid_en1 & ((\prif.pc_id [0])))

	.dataa(ifid_en),
	.datab(pc_0),
	.datac(prifpc_id_0),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_id1),
	.cout());
// synopsys translate_off
defparam \pc_id~1 .lut_mask = 16'hD8D8;
defparam \pc_id~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N4
cycloneive_lcell_comb \pc_id~2 (
// Equation(s):
// pc_id2 = (ifid_en1 & ((\Add2~0_combout ))) # (!ifid_en1 & (\prif.pc_id [3]))

	.dataa(gnd),
	.datab(ifid_en),
	.datac(prifpc_id_3),
	.datad(Add2),
	.cin(gnd),
	.combout(pc_id2),
	.cout());
// synopsys translate_off
defparam \pc_id~2 .lut_mask = 16'hFC30;
defparam \pc_id~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N16
cycloneive_lcell_comb \pc_id~3 (
// Equation(s):
// pc_id3 = (ifid_en1 & ((!pc_2))) # (!ifid_en1 & (\prif.pc_id [2]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifpc_id_2),
	.datad(pc_2),
	.cin(gnd),
	.combout(pc_id3),
	.cout());
// synopsys translate_off
defparam \pc_id~3 .lut_mask = 16'h50FA;
defparam \pc_id~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N22
cycloneive_lcell_comb \pc_id~4 (
// Equation(s):
// pc_id4 = (ifid_en1 & ((\Add2~4_combout ))) # (!ifid_en1 & (\prif.pc_id [5]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifpc_id_5),
	.datad(Add22),
	.cin(gnd),
	.combout(pc_id4),
	.cout());
// synopsys translate_off
defparam \pc_id~4 .lut_mask = 16'hFA50;
defparam \pc_id~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N6
cycloneive_lcell_comb \pc_id~5 (
// Equation(s):
// pc_id5 = (ifid_en1 & (\Add2~2_combout )) # (!ifid_en1 & ((\prif.pc_id [4])))

	.dataa(gnd),
	.datab(Add21),
	.datac(prifpc_id_4),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id5),
	.cout());
// synopsys translate_off
defparam \pc_id~5 .lut_mask = 16'hCCF0;
defparam \pc_id~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N4
cycloneive_lcell_comb \pc_id~6 (
// Equation(s):
// pc_id6 = (ifid_en1 & (\Add2~8_combout )) # (!ifid_en1 & ((\prif.pc_id [7])))

	.dataa(Add24),
	.datab(gnd),
	.datac(prifpc_id_7),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id6),
	.cout());
// synopsys translate_off
defparam \pc_id~6 .lut_mask = 16'hAAF0;
defparam \pc_id~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N30
cycloneive_lcell_comb \pc_id~7 (
// Equation(s):
// pc_id7 = (ifid_en1 & (\Add2~6_combout )) # (!ifid_en1 & ((\prif.pc_id [6])))

	.dataa(Add23),
	.datab(gnd),
	.datac(prifpc_id_6),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id7),
	.cout());
// synopsys translate_off
defparam \pc_id~7 .lut_mask = 16'hAAF0;
defparam \pc_id~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N20
cycloneive_lcell_comb \pc_id~8 (
// Equation(s):
// pc_id8 = (ifid_en1 & (\Add2~12_combout )) # (!ifid_en1 & ((\prif.pc_id [9])))

	.dataa(gnd),
	.datab(Add26),
	.datac(prifpc_id_9),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id8),
	.cout());
// synopsys translate_off
defparam \pc_id~8 .lut_mask = 16'hCCF0;
defparam \pc_id~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N18
cycloneive_lcell_comb \pc_id~9 (
// Equation(s):
// pc_id9 = (ifid_en1 & (\Add2~10_combout )) # (!ifid_en1 & ((\prif.pc_id [8])))

	.dataa(Add25),
	.datab(gnd),
	.datac(prifpc_id_8),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id9),
	.cout());
// synopsys translate_off
defparam \pc_id~9 .lut_mask = 16'hAAF0;
defparam \pc_id~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N0
cycloneive_lcell_comb \pc_id~10 (
// Equation(s):
// pc_id10 = (ifid_en1 & (\Add2~16_combout )) # (!ifid_en1 & ((\prif.pc_id [11])))

	.dataa(gnd),
	.datab(Add28),
	.datac(prifpc_id_11),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id10),
	.cout());
// synopsys translate_off
defparam \pc_id~10 .lut_mask = 16'hCCF0;
defparam \pc_id~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N12
cycloneive_lcell_comb \pc_id~11 (
// Equation(s):
// pc_id11 = (ifid_en1 & ((\Add2~14_combout ))) # (!ifid_en1 & (\prif.pc_id [10]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifpc_id_10),
	.datad(Add27),
	.cin(gnd),
	.combout(pc_id11),
	.cout());
// synopsys translate_off
defparam \pc_id~11 .lut_mask = 16'hFA50;
defparam \pc_id~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N28
cycloneive_lcell_comb \pc_id~12 (
// Equation(s):
// pc_id12 = (ifid_en1 & (\Add2~20_combout )) # (!ifid_en1 & ((\prif.pc_id [13])))

	.dataa(gnd),
	.datab(Add210),
	.datac(prifpc_id_13),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id12),
	.cout());
// synopsys translate_off
defparam \pc_id~12 .lut_mask = 16'hCCF0;
defparam \pc_id~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y33_N2
cycloneive_lcell_comb \pc_id~13 (
// Equation(s):
// pc_id13 = (ifid_en1 & (\Add2~18_combout )) # (!ifid_en1 & ((\prif.pc_id [12])))

	.dataa(Add29),
	.datab(gnd),
	.datac(prifpc_id_12),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id13),
	.cout());
// synopsys translate_off
defparam \pc_id~13 .lut_mask = 16'hAAF0;
defparam \pc_id~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N30
cycloneive_lcell_comb \pc_id~14 (
// Equation(s):
// pc_id14 = (ifid_en1 & ((\Add2~24_combout ))) # (!ifid_en1 & (\prif.pc_id [15]))

	.dataa(gnd),
	.datab(ifid_en),
	.datac(prifpc_id_15),
	.datad(Add212),
	.cin(gnd),
	.combout(pc_id14),
	.cout());
// synopsys translate_off
defparam \pc_id~14 .lut_mask = 16'hFC30;
defparam \pc_id~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N10
cycloneive_lcell_comb \pc_id~15 (
// Equation(s):
// pc_id15 = (ifid_en1 & (\Add2~22_combout )) # (!ifid_en1 & ((\prif.pc_id [14])))

	.dataa(Add211),
	.datab(gnd),
	.datac(prifpc_id_14),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id15),
	.cout());
// synopsys translate_off
defparam \pc_id~15 .lut_mask = 16'hAAF0;
defparam \pc_id~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y32_N30
cycloneive_lcell_comb \pc_id~16 (
// Equation(s):
// pc_id16 = (ifid_en1 & (\Add2~40_combout )) # (!ifid_en1 & ((\prif.pc_id [23])))

	.dataa(Add220),
	.datab(gnd),
	.datac(prifpc_id_23),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id16),
	.cout());
// synopsys translate_off
defparam \pc_id~16 .lut_mask = 16'hAAF0;
defparam \pc_id~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N12
cycloneive_lcell_comb \pc_id~17 (
// Equation(s):
// pc_id17 = (ifid_en1 & ((\Add2~38_combout ))) # (!ifid_en1 & (\prif.pc_id [22]))

	.dataa(gnd),
	.datab(ifid_en),
	.datac(prifpc_id_22),
	.datad(Add219),
	.cin(gnd),
	.combout(pc_id17),
	.cout());
// synopsys translate_off
defparam \pc_id~17 .lut_mask = 16'hFC30;
defparam \pc_id~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N24
cycloneive_lcell_comb \pc_id~18 (
// Equation(s):
// pc_id18 = (ifid_en1 & (\Add2~36_combout )) # (!ifid_en1 & ((\prif.pc_id [21])))

	.dataa(gnd),
	.datab(Add218),
	.datac(prifpc_id_21),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id18),
	.cout());
// synopsys translate_off
defparam \pc_id~18 .lut_mask = 16'hCCF0;
defparam \pc_id~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N2
cycloneive_lcell_comb \pc_id~19 (
// Equation(s):
// pc_id19 = (ifid_en1 & (\Add2~34_combout )) # (!ifid_en1 & ((\prif.pc_id [20])))

	.dataa(gnd),
	.datab(Add217),
	.datac(prifpc_id_20),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id19),
	.cout());
// synopsys translate_off
defparam \pc_id~19 .lut_mask = 16'hCCF0;
defparam \pc_id~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N16
cycloneive_lcell_comb \pc_id~20 (
// Equation(s):
// pc_id20 = (ifid_en1 & (\Add2~32_combout )) # (!ifid_en1 & ((\prif.pc_id [19])))

	.dataa(gnd),
	.datab(Add216),
	.datac(prifpc_id_19),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id20),
	.cout());
// synopsys translate_off
defparam \pc_id~20 .lut_mask = 16'hCCF0;
defparam \pc_id~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N14
cycloneive_lcell_comb \pc_id~21 (
// Equation(s):
// pc_id21 = (ifid_en1 & (\Add2~30_combout )) # (!ifid_en1 & ((\prif.pc_id [18])))

	.dataa(gnd),
	.datab(Add215),
	.datac(prifpc_id_18),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id21),
	.cout());
// synopsys translate_off
defparam \pc_id~21 .lut_mask = 16'hCCF0;
defparam \pc_id~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N0
cycloneive_lcell_comb \pc_id~22 (
// Equation(s):
// pc_id22 = (ifid_en1 & (\Add2~28_combout )) # (!ifid_en1 & ((\prif.pc_id [17])))

	.dataa(gnd),
	.datab(Add214),
	.datac(prifpc_id_17),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id22),
	.cout());
// synopsys translate_off
defparam \pc_id~22 .lut_mask = 16'hCCF0;
defparam \pc_id~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N22
cycloneive_lcell_comb \pc_id~23 (
// Equation(s):
// pc_id23 = (ifid_en1 & (\Add2~26_combout )) # (!ifid_en1 & ((\prif.pc_id [16])))

	.dataa(gnd),
	.datab(Add213),
	.datac(prifpc_id_16),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id23),
	.cout());
// synopsys translate_off
defparam \pc_id~23 .lut_mask = 16'hCCF0;
defparam \pc_id~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N12
cycloneive_lcell_comb \pc_id~24 (
// Equation(s):
// pc_id24 = (ifid_en1 & (\Add2~52_combout )) # (!ifid_en1 & ((\prif.pc_id [29])))

	.dataa(gnd),
	.datab(Add226),
	.datac(prifpc_id_29),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id24),
	.cout());
// synopsys translate_off
defparam \pc_id~24 .lut_mask = 16'hCCF0;
defparam \pc_id~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N18
cycloneive_lcell_comb \pc_id~25 (
// Equation(s):
// pc_id25 = (ifid_en1 & ((\Add2~50_combout ))) # (!ifid_en1 & (\prif.pc_id [28]))

	.dataa(gnd),
	.datab(ifid_en),
	.datac(prifpc_id_28),
	.datad(Add225),
	.cin(gnd),
	.combout(pc_id25),
	.cout());
// synopsys translate_off
defparam \pc_id~25 .lut_mask = 16'hFC30;
defparam \pc_id~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N0
cycloneive_lcell_comb \pc_id~26 (
// Equation(s):
// pc_id26 = (ifid_en1 & ((\Add2~48_combout ))) # (!ifid_en1 & (\prif.pc_id [27]))

	.dataa(gnd),
	.datab(ifid_en),
	.datac(prifpc_id_27),
	.datad(Add224),
	.cin(gnd),
	.combout(pc_id26),
	.cout());
// synopsys translate_off
defparam \pc_id~26 .lut_mask = 16'hFC30;
defparam \pc_id~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y32_N24
cycloneive_lcell_comb \pc_id~27 (
// Equation(s):
// pc_id27 = (ifid_en1 & (\Add2~46_combout )) # (!ifid_en1 & ((\prif.pc_id [26])))

	.dataa(Add223),
	.datab(gnd),
	.datac(prifpc_id_26),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id27),
	.cout());
// synopsys translate_off
defparam \pc_id~27 .lut_mask = 16'hAAF0;
defparam \pc_id~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X58_Y34_N26
cycloneive_lcell_comb \pc_id~28 (
// Equation(s):
// pc_id28 = (ifid_en1 & (\Add2~44_combout )) # (!ifid_en1 & ((\prif.pc_id [25])))

	.dataa(gnd),
	.datab(Add222),
	.datac(prifpc_id_25),
	.datad(ifid_en),
	.cin(gnd),
	.combout(pc_id28),
	.cout());
// synopsys translate_off
defparam \pc_id~28 .lut_mask = 16'hCCF0;
defparam \pc_id~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N14
cycloneive_lcell_comb \pc_id~29 (
// Equation(s):
// pc_id29 = (ifid_en1 & ((\Add2~42_combout ))) # (!ifid_en1 & (\prif.pc_id [24]))

	.dataa(ifid_en),
	.datab(gnd),
	.datac(prifpc_id_24),
	.datad(Add221),
	.cin(gnd),
	.combout(pc_id29),
	.cout());
// synopsys translate_off
defparam \pc_id~29 .lut_mask = 16'hFA50;
defparam \pc_id~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y34_N6
cycloneive_lcell_comb \pc_id~30 (
// Equation(s):
// pc_id30 = (ifid_en1 & ((\Add2~56_combout ))) # (!ifid_en1 & (\prif.pc_id [31]))

	.dataa(gnd),
	.datab(ifid_en),
	.datac(prifpc_id_31),
	.datad(Add228),
	.cin(gnd),
	.combout(pc_id30),
	.cout());
// synopsys translate_off
defparam \pc_id~30 .lut_mask = 16'hFC30;
defparam \pc_id~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N28
cycloneive_lcell_comb \pc_id~31 (
// Equation(s):
// pc_id31 = (ifid_en1 & (\Add2~54_combout )) # (!ifid_en1 & ((\prif.pc_id [30])))

	.dataa(ifid_en),
	.datab(Add227),
	.datac(prifpc_id_30),
	.datad(gnd),
	.cin(gnd),
	.combout(pc_id31),
	.cout());
// synopsys translate_off
defparam \pc_id~31 .lut_mask = 16'hD8D8;
defparam \pc_id~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y34_N30
cycloneive_lcell_comb \dataScr_ex~4 (
// Equation(s):
// dataScr_ex2 = (ccifiwait_0 & (((\prif.dataScr_ex [0])))) # (!ccifiwait_0 & (\prif.imemload_id [26] & ((Equal12))))

	.dataa(prifimemload_id_26),
	.datab(ccifiwait_0),
	.datac(prifdataScr_ex_0),
	.datad(Equal12),
	.cin(gnd),
	.combout(dataScr_ex2),
	.cout());
// synopsys translate_off
defparam \dataScr_ex~4 .lut_mask = 16'hE2C0;
defparam \dataScr_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N2
cycloneive_lcell_comb \ALUScr_ex~15 (
// Equation(s):
// ALUScr_ex3 = (!\prif.imemload_id [30] & ((\prif.imemload_id [26] & ((\ALUScr_ex~6_combout ))) # (!\prif.imemload_id [26] & (\ALUScr_ex~5_combout ))))

	.dataa(\ALUScr_ex~5_combout ),
	.datab(prifimemload_id_30),
	.datac(\ALUScr_ex~6_combout ),
	.datad(prifimemload_id_26),
	.cin(gnd),
	.combout(ALUScr_ex3),
	.cout());
// synopsys translate_off
defparam \ALUScr_ex~15 .lut_mask = 16'h3022;
defparam \ALUScr_ex~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N2
cycloneive_lcell_comb \zero_flag_mem~13 (
// Equation(s):
// zero_flag_mem = (exmem_en & (\zero_flag_mem~12_combout  & ((!\zero_flag_mem~2_combout )))) # (!exmem_en & (((\prif.zero_flag_mem~q ))))

	.dataa(exmem_en),
	.datab(\zero_flag_mem~12_combout ),
	.datac(prifzero_flag_mem),
	.datad(\zero_flag_mem~2_combout ),
	.cin(gnd),
	.combout(zero_flag_mem),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~13 .lut_mask = 16'h50D8;
defparam \zero_flag_mem~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N30
cycloneive_lcell_comb \ALUScr_ex~10 (
// Equation(s):
// \ALUScr_ex~10_combout  = ((\prif.imemload_id [27] & \prif.imemload_id [26])) # (!Equal20)

	.dataa(prifimemload_id_27),
	.datab(Equal20),
	.datac(gnd),
	.datad(prifimemload_id_26),
	.cin(gnd),
	.combout(\ALUScr_ex~10_combout ),
	.cout());
// synopsys translate_off
defparam \ALUScr_ex~10 .lut_mask = 16'hBB33;
defparam \ALUScr_ex~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N8
cycloneive_lcell_comb \ALUScr_ex~14 (
// Equation(s):
// \ALUScr_ex~14_combout  = ((Equal11 & (Equal0 & !\prif.imemload_id [3]))) # (!\ALUScr_ex~10_combout )

	.dataa(Equal11),
	.datab(Equal0),
	.datac(\ALUScr_ex~10_combout ),
	.datad(prifimemload_id_3),
	.cin(gnd),
	.combout(\ALUScr_ex~14_combout ),
	.cout());
// synopsys translate_off
defparam \ALUScr_ex~14 .lut_mask = 16'h0F8F;
defparam \ALUScr_ex~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N2
cycloneive_lcell_comb \ALUScr_ex~9 (
// Equation(s):
// \ALUScr_ex~9_combout  = ((\prif.imemload_id [26] & !\prif.imemload_id [28])) # (!Equal15)

	.dataa(gnd),
	.datab(Equal15),
	.datac(prifimemload_id_26),
	.datad(prifimemload_id_28),
	.cin(gnd),
	.combout(\ALUScr_ex~9_combout ),
	.cout());
// synopsys translate_off
defparam \ALUScr_ex~9 .lut_mask = 16'h33F3;
defparam \ALUScr_ex~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y30_N26
cycloneive_lcell_comb \regwrite_mem~0 (
// Equation(s):
// \regwrite_mem~0_combout  = (\prif.RegDest_ex [0] & (\prif.rd_ex [4] & (!\prif.RegDest_ex [1]))) # (!\prif.RegDest_ex [0] & (((\prif.RegDest_ex [1]) # (\prif.rt_ex [4]))))

	.dataa(prifrd_ex_4),
	.datab(prifRegDest_ex_0),
	.datac(prifRegDest_ex_1),
	.datad(prifrt_ex_4),
	.cin(gnd),
	.combout(\regwrite_mem~0_combout ),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~0 .lut_mask = 16'h3B38;
defparam \regwrite_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N26
cycloneive_lcell_comb \regwrite_mem~2 (
// Equation(s):
// \regwrite_mem~2_combout  = (\prif.RegDest_ex [0] & (\prif.rd_ex [0] & ((!\prif.RegDest_ex [1])))) # (!\prif.RegDest_ex [0] & (((\prif.rt_ex [0]) # (\prif.RegDest_ex [1]))))

	.dataa(prifRegDest_ex_0),
	.datab(prifrd_ex_0),
	.datac(prifrt_ex_0),
	.datad(prifRegDest_ex_1),
	.cin(gnd),
	.combout(\regwrite_mem~2_combout ),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~2 .lut_mask = 16'h55D8;
defparam \regwrite_mem~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X57_Y27_N6
cycloneive_lcell_comb \regwrite_mem~4 (
// Equation(s):
// \regwrite_mem~4_combout  = (\prif.RegDest_ex [1] & (((!\prif.RegDest_ex [0])))) # (!\prif.RegDest_ex [1] & ((\prif.RegDest_ex [0] & (\prif.rd_ex [1])) # (!\prif.RegDest_ex [0] & ((\prif.rt_ex [1])))))

	.dataa(prifrd_ex_1),
	.datab(prifRegDest_ex_1),
	.datac(prifRegDest_ex_0),
	.datad(prifrt_ex_1),
	.cin(gnd),
	.combout(\regwrite_mem~4_combout ),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~4 .lut_mask = 16'h2F2C;
defparam \regwrite_mem~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y33_N22
cycloneive_lcell_comb \regwrite_mem~6 (
// Equation(s):
// \regwrite_mem~6_combout  = (\prif.RegDest_ex [0] & (!\prif.RegDest_ex [1] & ((\prif.rd_ex [2])))) # (!\prif.RegDest_ex [0] & ((\prif.RegDest_ex [1]) # ((\prif.rt_ex [2]))))

	.dataa(prifRegDest_ex_0),
	.datab(prifRegDest_ex_1),
	.datac(prifrt_ex_2),
	.datad(prifrd_ex_2),
	.cin(gnd),
	.combout(\regwrite_mem~6_combout ),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~6 .lut_mask = 16'h7654;
defparam \regwrite_mem~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N12
cycloneive_lcell_comb \regwrite_mem~8 (
// Equation(s):
// \regwrite_mem~8_combout  = (\prif.RegDest_ex [1] & (((!\prif.RegDest_ex [0])))) # (!\prif.RegDest_ex [1] & ((\prif.RegDest_ex [0] & ((\prif.rd_ex [3]))) # (!\prif.RegDest_ex [0] & (\prif.rt_ex [3]))))

	.dataa(prifRegDest_ex_1),
	.datab(prifrt_ex_3),
	.datac(prifRegDest_ex_0),
	.datad(prifrd_ex_3),
	.cin(gnd),
	.combout(\regwrite_mem~8_combout ),
	.cout());
// synopsys translate_off
defparam \regwrite_mem~8 .lut_mask = 16'h5E0E;
defparam \regwrite_mem~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N16
cycloneive_lcell_comb \rdat2_ex~0 (
// Equation(s):
// \rdat2_ex~0_combout  = (\prif.imemload_id [20] & ((Mux62))) # (!\prif.imemload_id [20] & (Mux621))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux623),
	.datad(Mux622),
	.cin(gnd),
	.combout(\rdat2_ex~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~0 .lut_mask = 16'hFC30;
defparam \rdat2_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N18
cycloneive_lcell_comb \rdat1_ex~0 (
// Equation(s):
// \rdat1_ex~0_combout  = (\prif.imemload_id [25] & (Mux30)) # (!\prif.imemload_id [25] & ((Mux301)))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux30),
	.datad(Mux301),
	.cin(gnd),
	.combout(\rdat1_ex~0_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~0 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N2
cycloneive_lcell_comb \rdat2_ex~2 (
// Equation(s):
// \rdat2_ex~2_combout  = (\prif.imemload_id [20] & (Mux63)) # (!\prif.imemload_id [20] & ((Mux631)))

	.dataa(gnd),
	.datab(Mux632),
	.datac(Mux633),
	.datad(prifimemload_id_20),
	.cin(gnd),
	.combout(\rdat2_ex~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~2 .lut_mask = 16'hCCF0;
defparam \rdat2_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N16
cycloneive_lcell_comb \rdat1_ex~2 (
// Equation(s):
// \rdat1_ex~2_combout  = (\prif.imemload_id [25] & ((Mux31))) # (!\prif.imemload_id [25] & (Mux311))

	.dataa(Mux311),
	.datab(prifimemload_id_25),
	.datac(Mux31),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat1_ex~2_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~2 .lut_mask = 16'hE2E2;
defparam \rdat1_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y28_N16
cycloneive_lcell_comb \rdat2_ex~4 (
// Equation(s):
// \rdat2_ex~4_combout  = (\prif.imemload_id [20] & (Mux60)) # (!\prif.imemload_id [20] & ((Mux601)))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux60),
	.datad(Mux601),
	.cin(gnd),
	.combout(\rdat2_ex~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~4 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N28
cycloneive_lcell_comb \rdat2_ex~6 (
// Equation(s):
// \rdat2_ex~6_combout  = (\prif.imemload_id [20] & (Mux61)) # (!\prif.imemload_id [20] & ((Mux611)))

	.dataa(gnd),
	.datab(Mux611),
	.datac(Mux612),
	.datad(prifimemload_id_20),
	.cin(gnd),
	.combout(\rdat2_ex~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~6 .lut_mask = 16'hCCF0;
defparam \rdat2_ex~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N2
cycloneive_lcell_comb \rdat2_ex~8 (
// Equation(s):
// \rdat2_ex~8_combout  = (\prif.imemload_id [20] & ((Mux59))) # (!\prif.imemload_id [20] & (Mux591))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux591),
	.datad(Mux59),
	.cin(gnd),
	.combout(\rdat2_ex~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~8 .lut_mask = 16'hFC30;
defparam \rdat2_ex~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N14
cycloneive_lcell_comb \rdat2_ex~10 (
// Equation(s):
// \rdat2_ex~10_combout  = (\prif.imemload_id [20] & ((Mux32))) # (!\prif.imemload_id [20] & (Mux321))

	.dataa(prifimemload_id_20),
	.datab(gnd),
	.datac(Mux322),
	.datad(Mux321),
	.cin(gnd),
	.combout(\rdat2_ex~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~10 .lut_mask = 16'hFA50;
defparam \rdat2_ex~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N12
cycloneive_lcell_comb \rdat2_ex~12 (
// Equation(s):
// \rdat2_ex~12_combout  = (\prif.imemload_id [20] & ((Mux33))) # (!\prif.imemload_id [20] & (Mux331))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux332),
	.datad(Mux331),
	.cin(gnd),
	.combout(\rdat2_ex~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~12 .lut_mask = 16'hFC30;
defparam \rdat2_ex~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y27_N10
cycloneive_lcell_comb \rdat2_ex~14 (
// Equation(s):
// \rdat2_ex~14_combout  = (\prif.imemload_id [20] & ((Mux34))) # (!\prif.imemload_id [20] & (Mux341))

	.dataa(Mux342),
	.datab(prifimemload_id_20),
	.datac(Mux341),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat2_ex~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~14 .lut_mask = 16'hE2E2;
defparam \rdat2_ex~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N30
cycloneive_lcell_comb \rdat2_ex~16 (
// Equation(s):
// \rdat2_ex~16_combout  = (\prif.imemload_id [20] & ((Mux58))) # (!\prif.imemload_id [20] & (Mux581))

	.dataa(gnd),
	.datab(Mux581),
	.datac(prifimemload_id_20),
	.datad(Mux58),
	.cin(gnd),
	.combout(\rdat2_ex~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~16 .lut_mask = 16'hFC0C;
defparam \rdat2_ex~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N14
cycloneive_lcell_comb \rdat2_ex~18 (
// Equation(s):
// \rdat2_ex~18_combout  = (\prif.imemload_id [20] & (Mux48)) # (!\prif.imemload_id [20] & ((Mux481)))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux48),
	.datad(Mux481),
	.cin(gnd),
	.combout(\rdat2_ex~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~18 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N18
cycloneive_lcell_comb \rdat2_ex~20 (
// Equation(s):
// \rdat2_ex~20_combout  = (\prif.imemload_id [20] & ((Mux49))) # (!\prif.imemload_id [20] & (Mux491))

	.dataa(Mux491),
	.datab(Mux49),
	.datac(gnd),
	.datad(prifimemload_id_20),
	.cin(gnd),
	.combout(\rdat2_ex~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~20 .lut_mask = 16'hCCAA;
defparam \rdat2_ex~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N4
cycloneive_lcell_comb \rdat2_ex~22 (
// Equation(s):
// \rdat2_ex~22_combout  = (\prif.imemload_id [20] & ((Mux50))) # (!\prif.imemload_id [20] & (Mux501))

	.dataa(prifimemload_id_20),
	.datab(gnd),
	.datac(Mux501),
	.datad(Mux50),
	.cin(gnd),
	.combout(\rdat2_ex~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~22 .lut_mask = 16'hFA50;
defparam \rdat2_ex~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N6
cycloneive_lcell_comb \rdat2_ex~24 (
// Equation(s):
// \rdat2_ex~24_combout  = (\prif.imemload_id [20] & ((Mux51))) # (!\prif.imemload_id [20] & (Mux511))

	.dataa(prifimemload_id_20),
	.datab(gnd),
	.datac(Mux511),
	.datad(Mux51),
	.cin(gnd),
	.combout(\rdat2_ex~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~24 .lut_mask = 16'hFA50;
defparam \rdat2_ex~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N4
cycloneive_lcell_comb \rdat2_ex~26 (
// Equation(s):
// \rdat2_ex~26_combout  = (\prif.imemload_id [20] & ((Mux52))) # (!\prif.imemload_id [20] & (Mux521))

	.dataa(prifimemload_id_20),
	.datab(gnd),
	.datac(Mux521),
	.datad(Mux52),
	.cin(gnd),
	.combout(\rdat2_ex~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~26 .lut_mask = 16'hFA50;
defparam \rdat2_ex~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N0
cycloneive_lcell_comb \rdat2_ex~28 (
// Equation(s):
// \rdat2_ex~28_combout  = (\prif.imemload_id [20] & ((Mux53))) # (!\prif.imemload_id [20] & (Mux531))

	.dataa(gnd),
	.datab(Mux531),
	.datac(prifimemload_id_20),
	.datad(Mux53),
	.cin(gnd),
	.combout(\rdat2_ex~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~28 .lut_mask = 16'hFC0C;
defparam \rdat2_ex~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N30
cycloneive_lcell_comb \rdat2_ex~30 (
// Equation(s):
// \rdat2_ex~30_combout  = (\prif.imemload_id [20] & (Mux54)) # (!\prif.imemload_id [20] & ((Mux541)))

	.dataa(prifimemload_id_20),
	.datab(gnd),
	.datac(Mux54),
	.datad(Mux541),
	.cin(gnd),
	.combout(\rdat2_ex~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~30 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N16
cycloneive_lcell_comb \rdat2_ex~32 (
// Equation(s):
// \rdat2_ex~32_combout  = (\prif.imemload_id [20] & ((Mux57))) # (!\prif.imemload_id [20] & (Mux571))

	.dataa(prifimemload_id_20),
	.datab(Mux571),
	.datac(gnd),
	.datad(Mux57),
	.cin(gnd),
	.combout(\rdat2_ex~32_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~32 .lut_mask = 16'hEE44;
defparam \rdat2_ex~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N2
cycloneive_lcell_comb \rdat2_ex~34 (
// Equation(s):
// \rdat2_ex~34_combout  = (\prif.imemload_id [20] & ((Mux36))) # (!\prif.imemload_id [20] & (Mux361))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux362),
	.datad(Mux361),
	.cin(gnd),
	.combout(\rdat2_ex~34_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~34 .lut_mask = 16'hFC30;
defparam \rdat2_ex~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N8
cycloneive_lcell_comb \rdat2_ex~36 (
// Equation(s):
// \rdat2_ex~36_combout  = (\prif.imemload_id [20] & (Mux40)) # (!\prif.imemload_id [20] & ((Mux401)))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux401),
	.datad(Mux402),
	.cin(gnd),
	.combout(\rdat2_ex~36_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~36 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N10
cycloneive_lcell_comb \rdat2_ex~38 (
// Equation(s):
// \rdat2_ex~38_combout  = (\prif.imemload_id [20] & (Mux45)) # (!\prif.imemload_id [20] & ((Mux451)))

	.dataa(prifimemload_id_20),
	.datab(gnd),
	.datac(Mux451),
	.datad(Mux452),
	.cin(gnd),
	.combout(\rdat2_ex~38_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~38 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N0
cycloneive_lcell_comb \rdat2_ex~40 (
// Equation(s):
// \rdat2_ex~40_combout  = (\prif.imemload_id [20] & (Mux39)) # (!\prif.imemload_id [20] & ((Mux391)))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux391),
	.datad(Mux392),
	.cin(gnd),
	.combout(\rdat2_ex~40_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~40 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N18
cycloneive_lcell_comb \rdat2_ex~42 (
// Equation(s):
// \rdat2_ex~42_combout  = (\prif.imemload_id [20] & ((Mux47))) # (!\prif.imemload_id [20] & (Mux471))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux472),
	.datad(Mux471),
	.cin(gnd),
	.combout(\rdat2_ex~42_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~42 .lut_mask = 16'hFC30;
defparam \rdat2_ex~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N10
cycloneive_lcell_comb \rdat2_ex~44 (
// Equation(s):
// \rdat2_ex~44_combout  = (\prif.imemload_id [20] & ((Mux44))) # (!\prif.imemload_id [20] & (Mux441))

	.dataa(Mux442),
	.datab(Mux441),
	.datac(gnd),
	.datad(prifimemload_id_20),
	.cin(gnd),
	.combout(\rdat2_ex~44_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~44 .lut_mask = 16'hCCAA;
defparam \rdat2_ex~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N2
cycloneive_lcell_comb \rdat2_ex~46 (
// Equation(s):
// \rdat2_ex~46_combout  = (\prif.imemload_id [20] & ((Mux46))) # (!\prif.imemload_id [20] & (Mux461))

	.dataa(prifimemload_id_20),
	.datab(Mux462),
	.datac(gnd),
	.datad(Mux461),
	.cin(gnd),
	.combout(\rdat2_ex~46_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~46 .lut_mask = 16'hEE44;
defparam \rdat2_ex~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N6
cycloneive_lcell_comb \rdat2_ex~48 (
// Equation(s):
// \rdat2_ex~48_combout  = (\prif.imemload_id [20] & ((Mux42))) # (!\prif.imemload_id [20] & (Mux421))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux422),
	.datad(Mux421),
	.cin(gnd),
	.combout(\rdat2_ex~48_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~48 .lut_mask = 16'hFC30;
defparam \rdat2_ex~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N6
cycloneive_lcell_comb \rdat2_ex~50 (
// Equation(s):
// \rdat2_ex~50_combout  = (\prif.imemload_id [20] & (Mux43)) # (!\prif.imemload_id [20] & ((Mux431)))

	.dataa(prifimemload_id_20),
	.datab(gnd),
	.datac(Mux431),
	.datad(Mux432),
	.cin(gnd),
	.combout(\rdat2_ex~50_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~50 .lut_mask = 16'hF5A0;
defparam \rdat2_ex~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N0
cycloneive_lcell_comb \rdat2_ex~52 (
// Equation(s):
// \rdat2_ex~52_combout  = (\prif.imemload_id [20] & ((Mux35))) # (!\prif.imemload_id [20] & (Mux351))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux352),
	.datad(Mux351),
	.cin(gnd),
	.combout(\rdat2_ex~52_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~52 .lut_mask = 16'hFC30;
defparam \rdat2_ex~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N2
cycloneive_lcell_comb \rdat2_ex~54 (
// Equation(s):
// \rdat2_ex~54_combout  = (\prif.imemload_id [20] & (Mux37)) # (!\prif.imemload_id [20] & ((Mux371)))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux371),
	.datad(Mux372),
	.cin(gnd),
	.combout(\rdat2_ex~54_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~54 .lut_mask = 16'hF3C0;
defparam \rdat2_ex~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N24
cycloneive_lcell_comb \rdat2_ex~56 (
// Equation(s):
// \rdat2_ex~56_combout  = (\prif.imemload_id [20] & ((Mux55))) # (!\prif.imemload_id [20] & (Mux551))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux551),
	.datad(Mux55),
	.cin(gnd),
	.combout(\rdat2_ex~56_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~56 .lut_mask = 16'hFC30;
defparam \rdat2_ex~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N20
cycloneive_lcell_comb \rdat2_ex~58 (
// Equation(s):
// \rdat2_ex~58_combout  = (\prif.imemload_id [20] & ((Mux56))) # (!\prif.imemload_id [20] & (Mux561))

	.dataa(prifimemload_id_20),
	.datab(gnd),
	.datac(Mux561),
	.datad(Mux56),
	.cin(gnd),
	.combout(\rdat2_ex~58_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~58 .lut_mask = 16'hFA50;
defparam \rdat2_ex~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N6
cycloneive_lcell_comb \rdat2_ex~60 (
// Equation(s):
// \rdat2_ex~60_combout  = (\prif.imemload_id [20] & ((Mux41))) # (!\prif.imemload_id [20] & (Mux411))

	.dataa(gnd),
	.datab(prifimemload_id_20),
	.datac(Mux412),
	.datad(Mux411),
	.cin(gnd),
	.combout(\rdat2_ex~60_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~60 .lut_mask = 16'hFC30;
defparam \rdat2_ex~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y28_N0
cycloneive_lcell_comb \rdat2_ex~62 (
// Equation(s):
// \rdat2_ex~62_combout  = (\prif.imemload_id [20] & ((Mux38))) # (!\prif.imemload_id [20] & (Mux381))

	.dataa(prifimemload_id_20),
	.datab(Mux382),
	.datac(gnd),
	.datad(Mux381),
	.cin(gnd),
	.combout(\rdat2_ex~62_combout ),
	.cout());
// synopsys translate_off
defparam \rdat2_ex~62 .lut_mask = 16'hEE44;
defparam \rdat2_ex~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N18
cycloneive_lcell_comb \ALUOP_ex~1 (
// Equation(s):
// \ALUOP_ex~1_combout  = ((Equal4 & Equal11)) # (!\ALUScr_ex~10_combout )

	.dataa(\ALUScr_ex~10_combout ),
	.datab(Equal4),
	.datac(Equal11),
	.datad(gnd),
	.cin(gnd),
	.combout(\ALUOP_ex~1_combout ),
	.cout());
// synopsys translate_off
defparam \ALUOP_ex~1 .lut_mask = 16'hD5D5;
defparam \ALUOP_ex~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y25_N2
cycloneive_lcell_comb \rdat1_ex~4 (
// Equation(s):
// \rdat1_ex~4_combout  = (\prif.imemload_id [25] & ((Mux29))) # (!\prif.imemload_id [25] & (Mux291))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux291),
	.datad(Mux29),
	.cin(gnd),
	.combout(\rdat1_ex~4_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~4 .lut_mask = 16'hFC30;
defparam \rdat1_ex~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N0
cycloneive_lcell_comb \rdat1_ex~6 (
// Equation(s):
// \rdat1_ex~6_combout  = (\prif.imemload_id [25] & ((Mux27))) # (!\prif.imemload_id [25] & (Mux271))

	.dataa(Mux271),
	.datab(gnd),
	.datac(prifimemload_id_25),
	.datad(Mux27),
	.cin(gnd),
	.combout(\rdat1_ex~6_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~6 .lut_mask = 16'hFA0A;
defparam \rdat1_ex~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N12
cycloneive_lcell_comb \rdat1_ex~8 (
// Equation(s):
// \rdat1_ex~8_combout  = (\prif.imemload_id [25] & ((Mux28))) # (!\prif.imemload_id [25] & (Mux281))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux281),
	.datad(Mux28),
	.cin(gnd),
	.combout(\rdat1_ex~8_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~8 .lut_mask = 16'hFC30;
defparam \rdat1_ex~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N20
cycloneive_lcell_comb \rdat1_ex~10 (
// Equation(s):
// \rdat1_ex~10_combout  = (\prif.imemload_id [25] & ((Mux23))) # (!\prif.imemload_id [25] & (Mux231))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux231),
	.datad(Mux23),
	.cin(gnd),
	.combout(\rdat1_ex~10_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~10 .lut_mask = 16'hFC30;
defparam \rdat1_ex~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N14
cycloneive_lcell_comb \rdat1_ex~12 (
// Equation(s):
// \rdat1_ex~12_combout  = (\prif.imemload_id [25] & ((Mux24))) # (!\prif.imemload_id [25] & (Mux241))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux241),
	.datad(Mux24),
	.cin(gnd),
	.combout(\rdat1_ex~12_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~12 .lut_mask = 16'hFC30;
defparam \rdat1_ex~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N18
cycloneive_lcell_comb \rdat1_ex~14 (
// Equation(s):
// \rdat1_ex~14_combout  = (\prif.imemload_id [25] & ((Mux25))) # (!\prif.imemload_id [25] & (Mux251))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux251),
	.datad(Mux25),
	.cin(gnd),
	.combout(\rdat1_ex~14_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~14 .lut_mask = 16'hFC30;
defparam \rdat1_ex~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N18
cycloneive_lcell_comb \rdat1_ex~16 (
// Equation(s):
// \rdat1_ex~16_combout  = (\prif.imemload_id [25] & (Mux26)) # (!\prif.imemload_id [25] & ((Mux261)))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux26),
	.datad(Mux261),
	.cin(gnd),
	.combout(\rdat1_ex~16_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~16 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N6
cycloneive_lcell_comb \rdat1_ex~18 (
// Equation(s):
// \rdat1_ex~18_combout  = (\prif.imemload_id [25] & ((Mux15))) # (!\prif.imemload_id [25] & (Mux1510))

	.dataa(prifimemload_id_25),
	.datab(Mux151),
	.datac(gnd),
	.datad(Mux15),
	.cin(gnd),
	.combout(\rdat1_ex~18_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~18 .lut_mask = 16'hEE44;
defparam \rdat1_ex~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N12
cycloneive_lcell_comb \rdat1_ex~20 (
// Equation(s):
// \rdat1_ex~20_combout  = (\prif.imemload_id [25] & ((Mux16))) # (!\prif.imemload_id [25] & (Mux165))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux161),
	.datad(Mux16),
	.cin(gnd),
	.combout(\rdat1_ex~20_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~20 .lut_mask = 16'hFC30;
defparam \rdat1_ex~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N2
cycloneive_lcell_comb \rdat1_ex~22 (
// Equation(s):
// \rdat1_ex~22_combout  = (\prif.imemload_id [25] & (Mux17)) # (!\prif.imemload_id [25] & ((Mux171)))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux17),
	.datad(Mux171),
	.cin(gnd),
	.combout(\rdat1_ex~22_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~22 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N24
cycloneive_lcell_comb \rdat1_ex~24 (
// Equation(s):
// \rdat1_ex~24_combout  = (\prif.imemload_id [25] & ((Mux18))) # (!\prif.imemload_id [25] & (Mux181))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux181),
	.datad(Mux18),
	.cin(gnd),
	.combout(\rdat1_ex~24_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~24 .lut_mask = 16'hFC30;
defparam \rdat1_ex~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N12
cycloneive_lcell_comb \rdat1_ex~26 (
// Equation(s):
// \rdat1_ex~26_combout  = (\prif.imemload_id [25] & (Mux20)) # (!\prif.imemload_id [25] & ((Mux201)))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux20),
	.datad(Mux201),
	.cin(gnd),
	.combout(\rdat1_ex~26_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~26 .lut_mask = 16'hF3C0;
defparam \rdat1_ex~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N18
cycloneive_lcell_comb \rdat1_ex~28 (
// Equation(s):
// \rdat1_ex~28_combout  = (\prif.imemload_id [25] & (Mux19)) # (!\prif.imemload_id [25] & ((Mux191)))

	.dataa(Mux19),
	.datab(Mux191),
	.datac(prifimemload_id_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat1_ex~28_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~28 .lut_mask = 16'hACAC;
defparam \rdat1_ex~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N24
cycloneive_lcell_comb \rdat1_ex~30 (
// Equation(s):
// \rdat1_ex~30_combout  = (\prif.imemload_id [25] & ((Mux21))) # (!\prif.imemload_id [25] & (Mux211))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux211),
	.datad(Mux21),
	.cin(gnd),
	.combout(\rdat1_ex~30_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~30 .lut_mask = 16'hFC30;
defparam \rdat1_ex~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N30
cycloneive_lcell_comb \rdat1_ex~32 (
// Equation(s):
// \rdat1_ex~32_combout  = (\prif.imemload_id [25] & ((Mux22))) # (!\prif.imemload_id [25] & (Mux221))

	.dataa(gnd),
	.datab(Mux221),
	.datac(prifimemload_id_25),
	.datad(Mux22),
	.cin(gnd),
	.combout(\rdat1_ex~32_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~32 .lut_mask = 16'hFC0C;
defparam \rdat1_ex~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N6
cycloneive_lcell_comb \rdat1_ex~34 (
// Equation(s):
// \rdat1_ex~34_combout  = (\prif.imemload_id [25] & ((Mux13))) # (!\prif.imemload_id [25] & (Mux131))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux131),
	.datad(Mux13),
	.cin(gnd),
	.combout(\rdat1_ex~34_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~34 .lut_mask = 16'hFC30;
defparam \rdat1_ex~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N18
cycloneive_lcell_comb \rdat1_ex~36 (
// Equation(s):
// \rdat1_ex~36_combout  = (\prif.imemload_id [25] & ((Mux14))) # (!\prif.imemload_id [25] & (Mux1410))

	.dataa(Mux141),
	.datab(Mux14),
	.datac(gnd),
	.datad(prifimemload_id_25),
	.cin(gnd),
	.combout(\rdat1_ex~36_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~36 .lut_mask = 16'hCCAA;
defparam \rdat1_ex~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N16
cycloneive_lcell_comb \rdat1_ex~38 (
// Equation(s):
// \rdat1_ex~38_combout  = (\prif.imemload_id [25] & ((Mux11))) # (!\prif.imemload_id [25] & (Mux111))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux111),
	.datad(Mux11),
	.cin(gnd),
	.combout(\rdat1_ex~38_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~38 .lut_mask = 16'hFC30;
defparam \rdat1_ex~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N26
cycloneive_lcell_comb \rdat1_ex~40 (
// Equation(s):
// \rdat1_ex~40_combout  = (\prif.imemload_id [25] & ((Mux12))) # (!\prif.imemload_id [25] & (Mux121))

	.dataa(prifimemload_id_25),
	.datab(gnd),
	.datac(Mux121),
	.datad(Mux12),
	.cin(gnd),
	.combout(\rdat1_ex~40_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~40 .lut_mask = 16'hFA50;
defparam \rdat1_ex~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N24
cycloneive_lcell_comb \rdat1_ex~42 (
// Equation(s):
// \rdat1_ex~42_combout  = (\prif.imemload_id [25] & (Mux9)) # (!\prif.imemload_id [25] & ((Mux91)))

	.dataa(Mux9),
	.datab(gnd),
	.datac(Mux91),
	.datad(prifimemload_id_25),
	.cin(gnd),
	.combout(\rdat1_ex~42_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~42 .lut_mask = 16'hAAF0;
defparam \rdat1_ex~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N28
cycloneive_lcell_comb \rdat1_ex~44 (
// Equation(s):
// \rdat1_ex~44_combout  = (\prif.imemload_id [25] & ((Mux10))) # (!\prif.imemload_id [25] & (Mux101))

	.dataa(Mux101),
	.datab(Mux10),
	.datac(prifimemload_id_25),
	.datad(gnd),
	.cin(gnd),
	.combout(\rdat1_ex~44_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~44 .lut_mask = 16'hCACA;
defparam \rdat1_ex~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N20
cycloneive_lcell_comb \rdat1_ex~46 (
// Equation(s):
// \rdat1_ex~46_combout  = (\prif.imemload_id [25] & (Mux7)) # (!\prif.imemload_id [25] & ((Mux71)))

	.dataa(prifimemload_id_25),
	.datab(gnd),
	.datac(Mux7),
	.datad(Mux71),
	.cin(gnd),
	.combout(\rdat1_ex~46_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~46 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N16
cycloneive_lcell_comb \rdat1_ex~48 (
// Equation(s):
// \rdat1_ex~48_combout  = (\prif.imemload_id [25] & (Mux8)) # (!\prif.imemload_id [25] & ((Mux81)))

	.dataa(Mux8),
	.datab(gnd),
	.datac(prifimemload_id_25),
	.datad(Mux81),
	.cin(gnd),
	.combout(\rdat1_ex~48_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~48 .lut_mask = 16'hAFA0;
defparam \rdat1_ex~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N18
cycloneive_lcell_comb \rdat1_ex~50 (
// Equation(s):
// \rdat1_ex~50_combout  = (\prif.imemload_id [25] & (Mux0)) # (!\prif.imemload_id [25] & ((Mux01)))

	.dataa(prifimemload_id_25),
	.datab(gnd),
	.datac(Mux0),
	.datad(Mux01),
	.cin(gnd),
	.combout(\rdat1_ex~50_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~50 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~50 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N24
cycloneive_lcell_comb \rdat1_ex~52 (
// Equation(s):
// \rdat1_ex~52_combout  = (\prif.imemload_id [25] & ((Mux1))) # (!\prif.imemload_id [25] & (Mux110))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux110),
	.datad(Mux1),
	.cin(gnd),
	.combout(\rdat1_ex~52_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~52 .lut_mask = 16'hFC30;
defparam \rdat1_ex~52 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N14
cycloneive_lcell_comb \rdat1_ex~54 (
// Equation(s):
// \rdat1_ex~54_combout  = (\prif.imemload_id [25] & ((Mux2))) # (!\prif.imemload_id [25] & (Mux210))

	.dataa(gnd),
	.datab(prifimemload_id_25),
	.datac(Mux210),
	.datad(Mux2),
	.cin(gnd),
	.combout(\rdat1_ex~54_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~54 .lut_mask = 16'hFC30;
defparam \rdat1_ex~54 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N26
cycloneive_lcell_comb \rdat1_ex~56 (
// Equation(s):
// \rdat1_ex~56_combout  = (\prif.imemload_id [25] & (Mux5)) # (!\prif.imemload_id [25] & ((Mux510)))

	.dataa(Mux5),
	.datab(prifimemload_id_25),
	.datac(gnd),
	.datad(Mux510),
	.cin(gnd),
	.combout(\rdat1_ex~56_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~56 .lut_mask = 16'hBB88;
defparam \rdat1_ex~56 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N28
cycloneive_lcell_comb \rdat1_ex~58 (
// Equation(s):
// \rdat1_ex~58_combout  = (\prif.imemload_id [25] & (Mux6)) # (!\prif.imemload_id [25] & ((Mux64)))

	.dataa(prifimemload_id_25),
	.datab(gnd),
	.datac(Mux6),
	.datad(Mux64),
	.cin(gnd),
	.combout(\rdat1_ex~58_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~58 .lut_mask = 16'hF5A0;
defparam \rdat1_ex~58 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N6
cycloneive_lcell_comb \rdat1_ex~60 (
// Equation(s):
// \rdat1_ex~60_combout  = (\prif.imemload_id [25] & ((Mux3))) # (!\prif.imemload_id [25] & (Mux310))

	.dataa(prifimemload_id_25),
	.datab(gnd),
	.datac(Mux310),
	.datad(Mux3),
	.cin(gnd),
	.combout(\rdat1_ex~60_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~60 .lut_mask = 16'hFA50;
defparam \rdat1_ex~60 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N2
cycloneive_lcell_comb \rdat1_ex~62 (
// Equation(s):
// \rdat1_ex~62_combout  = (\prif.imemload_id [25] & (Mux4)) # (!\prif.imemload_id [25] & ((Mux410)))

	.dataa(Mux4),
	.datab(prifimemload_id_25),
	.datac(gnd),
	.datad(Mux410),
	.cin(gnd),
	.combout(\rdat1_ex~62_combout ),
	.cout());
// synopsys translate_off
defparam \rdat1_ex~62 .lut_mask = 16'hBB88;
defparam \rdat1_ex~62 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N16
cycloneive_lcell_comb \PCScr_ex~2 (
// Equation(s):
// \PCScr_ex~2_combout  = (\prif.imemload_id [31]) # (!Equal12)

	.dataa(prifimemload_id_31),
	.datab(gnd),
	.datac(gnd),
	.datad(Equal12),
	.cin(gnd),
	.combout(\PCScr_ex~2_combout ),
	.cout());
// synopsys translate_off
defparam \PCScr_ex~2 .lut_mask = 16'hAAFF;
defparam \PCScr_ex~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y32_N6
cycloneive_lcell_comb \PCScr_ex~5 (
// Equation(s):
// \PCScr_ex~5_combout  = (Equal10 & (Equal12 & ((!\prif.imemload_id [31])))) # (!Equal10 & ((Equal11) # ((Equal12 & !\prif.imemload_id [31]))))

	.dataa(Equal10),
	.datab(Equal12),
	.datac(Equal11),
	.datad(prifimemload_id_31),
	.cin(gnd),
	.combout(\PCScr_ex~5_combout ),
	.cout());
// synopsys translate_off
defparam \PCScr_ex~5 .lut_mask = 16'h50DC;
defparam \PCScr_ex~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N22
cycloneive_lcell_comb \ALUScr_ex~5 (
// Equation(s):
// \ALUScr_ex~5_combout  = (!\prif.imemload_id [31] & ((\prif.imemload_id [29]) # (!\prif.imemload_id [27])))

	.dataa(prifimemload_id_27),
	.datab(prifimemload_id_31),
	.datac(prifimemload_id_29),
	.datad(gnd),
	.cin(gnd),
	.combout(\ALUScr_ex~5_combout ),
	.cout());
// synopsys translate_off
defparam \ALUScr_ex~5 .lut_mask = 16'h3131;
defparam \ALUScr_ex~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y33_N4
cycloneive_lcell_comb \ALUScr_ex~6 (
// Equation(s):
// \ALUScr_ex~6_combout  = (\prif.imemload_id [28] & (((!\prif.imemload_id [31] & !\prif.imemload_id [27])))) # (!\prif.imemload_id [28] & ((\prif.imemload_id [31] & ((\prif.imemload_id [27]))) # (!\prif.imemload_id [31] & (\prif.imemload_id [29]))))

	.dataa(prifimemload_id_29),
	.datab(prifimemload_id_28),
	.datac(prifimemload_id_31),
	.datad(prifimemload_id_27),
	.cin(gnd),
	.combout(\ALUScr_ex~6_combout ),
	.cout());
// synopsys translate_off
defparam \ALUScr_ex~6 .lut_mask = 16'h320E;
defparam \ALUScr_ex~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y21_N10
cycloneive_lcell_comb \zero_flag_mem~0 (
// Equation(s):
// \zero_flag_mem~0_combout  = (!aluifportOut_3 & (!aluifportOut_21 & ((!aluifportOut_2) # (!aluifportOut_31))))

	.dataa(aluifportOut_31),
	.datab(aluifportOut_2),
	.datac(aluifportOut_3),
	.datad(aluifportOut_21),
	.cin(gnd),
	.combout(\zero_flag_mem~0_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~0 .lut_mask = 16'h0007;
defparam \zero_flag_mem~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y25_N14
cycloneive_lcell_comb \zero_flag_mem~6 (
// Equation(s):
// \zero_flag_mem~6_combout  = ((!aluifportOut_13 & (!aluifportOut_14 & !aluifportOut_15))) # (!\prif.ALUOP_ex [3])

	.dataa(aluifportOut_13),
	.datab(aluifportOut_14),
	.datac(prifALUOP_ex_3),
	.datad(aluifportOut_15),
	.cin(gnd),
	.combout(\zero_flag_mem~6_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~6 .lut_mask = 16'h0F1F;
defparam \zero_flag_mem~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N8
cycloneive_lcell_comb \zero_flag_mem~9 (
// Equation(s):
// \zero_flag_mem~9_combout  = ((!aluifportOut_20 & (!aluifportOut_211 & !aluifportOut_22))) # (!\prif.ALUOP_ex [3])

	.dataa(prifALUOP_ex_3),
	.datab(aluifportOut_20),
	.datac(aluifportOut_211),
	.datad(aluifportOut_22),
	.cin(gnd),
	.combout(\zero_flag_mem~9_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~9 .lut_mask = 16'h5557;
defparam \zero_flag_mem~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N12
cycloneive_lcell_comb \zero_flag_mem~7 (
// Equation(s):
// \zero_flag_mem~7_combout  = ((!aluifportOut_11 & (!aluifportOut_10 & !aluifportOut_9))) # (!\prif.ALUOP_ex [3])

	.dataa(prifALUOP_ex_3),
	.datab(aluifportOut_11),
	.datac(aluifportOut_10),
	.datad(aluifportOut_9),
	.cin(gnd),
	.combout(\zero_flag_mem~7_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~7 .lut_mask = 16'h5557;
defparam \zero_flag_mem~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N6
cycloneive_lcell_comb \zero_flag_mem~10 (
// Equation(s):
// \zero_flag_mem~10_combout  = (\zero_flag_mem~8_combout  & (\zero_flag_mem~6_combout  & (\zero_flag_mem~9_combout  & \zero_flag_mem~7_combout )))

	.dataa(\zero_flag_mem~8_combout ),
	.datab(\zero_flag_mem~6_combout ),
	.datac(\zero_flag_mem~9_combout ),
	.datad(\zero_flag_mem~7_combout ),
	.cin(gnd),
	.combout(\zero_flag_mem~10_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~10 .lut_mask = 16'h8000;
defparam \zero_flag_mem~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N28
cycloneive_lcell_comb \zero_flag_mem~11 (
// Equation(s):
// \zero_flag_mem~11_combout  = (\zero_flag_mem~5_combout  & (!aluifportOut_29 & (!aluifportOut_28 & \zero_flag_mem~10_combout )))

	.dataa(\zero_flag_mem~5_combout ),
	.datab(aluifportOut_29),
	.datac(aluifportOut_28),
	.datad(\zero_flag_mem~10_combout ),
	.cin(gnd),
	.combout(\zero_flag_mem~11_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~11 .lut_mask = 16'h0200;
defparam \zero_flag_mem~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N14
cycloneive_lcell_comb \zero_flag_mem~12 (
// Equation(s):
// \zero_flag_mem~12_combout  = (\zero_flag_mem~0_combout  & (!aluifportOut_1 & (!aluifportOut_0 & \zero_flag_mem~11_combout )))

	.dataa(\zero_flag_mem~0_combout ),
	.datab(aluifportOut_1),
	.datac(aluifportOut_0),
	.datad(\zero_flag_mem~11_combout ),
	.cin(gnd),
	.combout(\zero_flag_mem~12_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~12 .lut_mask = 16'h0200;
defparam \zero_flag_mem~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N10
cycloneive_lcell_comb \zero_flag_mem~1 (
// Equation(s):
// \zero_flag_mem~1_combout  = (aluifportOut_30) # ((aluifportOut_16) # ((aluifportOut_17) # (aluifportOut_19)))

	.dataa(aluifportOut_30),
	.datab(aluifportOut_16),
	.datac(aluifportOut_17),
	.datad(aluifportOut_19),
	.cin(gnd),
	.combout(\zero_flag_mem~1_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~1 .lut_mask = 16'hFFFE;
defparam \zero_flag_mem~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y25_N0
cycloneive_lcell_comb \zero_flag_mem~2 (
// Equation(s):
// \zero_flag_mem~2_combout  = (\prif.ALUOP_ex [3] & ((aluifneg_flag) # ((aluifportOut_18) # (\zero_flag_mem~1_combout ))))

	.dataa(prifALUOP_ex_3),
	.datab(aluifneg_flag),
	.datac(aluifportOut_18),
	.datad(\zero_flag_mem~1_combout ),
	.cin(gnd),
	.combout(\zero_flag_mem~2_combout ),
	.cout());
// synopsys translate_off
defparam \zero_flag_mem~2 .lut_mask = 16'hAAA8;
defparam \zero_flag_mem~2 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module register_file (
	prifimemload_id_17,
	prifimemload_id_16,
	prifimemload_id_19,
	prifimemload_id_18,
	prifimemload_id_22,
	prifimemload_id_21,
	prifimemload_id_24,
	prifimemload_id_23,
	prifRegwen_wb,
	prifregwrite_wb_2,
	prifregwrite_wb_0,
	prifregwrite_wb_1,
	prifregwrite_wb_4,
	prifregwrite_wb_3,
	Equal8,
	Mux163,
	Mux164,
	Mux161,
	Mux162,
	Mux160,
	Mux133,
	Mux134,
	Mux135,
	Mux159,
	Mux149,
	Mux150,
	Mux151,
	Mux152,
	Mux153,
	Mux154,
	Mux155,
	Mux158,
	Mux137,
	Mux141,
	Mux146,
	Mux140,
	Mux148,
	Mux145,
	Mux147,
	Mux143,
	Mux144,
	Mux136,
	Mux138,
	Mux156,
	Mux157,
	Mux142,
	Mux139,
	Mux62,
	Mux621,
	Mux30,
	Mux301,
	Mux63,
	Mux631,
	Mux31,
	Mux311,
	Mux60,
	Mux601,
	Mux61,
	Mux611,
	Mux59,
	Mux591,
	Mux32,
	Mux321,
	Mux33,
	Mux331,
	Mux34,
	Mux341,
	Mux58,
	Mux581,
	Mux48,
	Mux481,
	Mux49,
	Mux491,
	Mux50,
	Mux501,
	Mux51,
	Mux511,
	Mux52,
	Mux521,
	Mux53,
	Mux531,
	Mux54,
	Mux541,
	Mux57,
	Mux571,
	Mux36,
	Mux361,
	Mux40,
	Mux401,
	Mux45,
	Mux451,
	Mux39,
	Mux391,
	Mux47,
	Mux471,
	Mux44,
	Mux441,
	Mux46,
	Mux461,
	Mux42,
	Mux421,
	Mux43,
	Mux431,
	Mux35,
	Mux351,
	Mux37,
	Mux371,
	Mux55,
	Mux551,
	Mux56,
	Mux561,
	Mux41,
	Mux411,
	Mux38,
	Mux381,
	Mux29,
	Mux291,
	Mux27,
	Mux271,
	Mux28,
	Mux281,
	Mux23,
	Mux231,
	Mux24,
	Mux241,
	Mux25,
	Mux251,
	Mux26,
	Mux261,
	Mux15,
	Mux1510,
	Mux16,
	Mux165,
	Mux17,
	Mux171,
	Mux18,
	Mux181,
	Mux20,
	Mux201,
	Mux19,
	Mux191,
	Mux21,
	Mux211,
	Mux22,
	Mux221,
	Mux13,
	Mux131,
	Mux14,
	Mux1410,
	Mux11,
	Mux111,
	Mux12,
	Mux121,
	Mux9,
	Mux91,
	Mux10,
	Mux101,
	Mux7,
	Mux71,
	Mux8,
	Mux81,
	Mux0,
	Mux01,
	Mux1,
	Mux110,
	Mux2,
	Mux210,
	Mux5,
	Mux510,
	Mux6,
	Mux64,
	Mux3,
	Mux310,
	Mux4,
	Mux410,
	CLK,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	prifimemload_id_17;
input 	prifimemload_id_16;
input 	prifimemload_id_19;
input 	prifimemload_id_18;
input 	prifimemload_id_22;
input 	prifimemload_id_21;
input 	prifimemload_id_24;
input 	prifimemload_id_23;
input 	prifRegwen_wb;
input 	prifregwrite_wb_2;
input 	prifregwrite_wb_0;
input 	prifregwrite_wb_1;
input 	prifregwrite_wb_4;
input 	prifregwrite_wb_3;
input 	Equal8;
input 	Mux163;
input 	Mux164;
input 	Mux161;
input 	Mux162;
input 	Mux160;
input 	Mux133;
input 	Mux134;
input 	Mux135;
input 	Mux159;
input 	Mux149;
input 	Mux150;
input 	Mux151;
input 	Mux152;
input 	Mux153;
input 	Mux154;
input 	Mux155;
input 	Mux158;
input 	Mux137;
input 	Mux141;
input 	Mux146;
input 	Mux140;
input 	Mux148;
input 	Mux145;
input 	Mux147;
input 	Mux143;
input 	Mux144;
input 	Mux136;
input 	Mux138;
input 	Mux156;
input 	Mux157;
input 	Mux142;
input 	Mux139;
output 	Mux62;
output 	Mux621;
output 	Mux30;
output 	Mux301;
output 	Mux63;
output 	Mux631;
output 	Mux31;
output 	Mux311;
output 	Mux60;
output 	Mux601;
output 	Mux61;
output 	Mux611;
output 	Mux59;
output 	Mux591;
output 	Mux32;
output 	Mux321;
output 	Mux33;
output 	Mux331;
output 	Mux34;
output 	Mux341;
output 	Mux58;
output 	Mux581;
output 	Mux48;
output 	Mux481;
output 	Mux49;
output 	Mux491;
output 	Mux50;
output 	Mux501;
output 	Mux51;
output 	Mux511;
output 	Mux52;
output 	Mux521;
output 	Mux53;
output 	Mux531;
output 	Mux54;
output 	Mux541;
output 	Mux57;
output 	Mux571;
output 	Mux36;
output 	Mux361;
output 	Mux40;
output 	Mux401;
output 	Mux45;
output 	Mux451;
output 	Mux39;
output 	Mux391;
output 	Mux47;
output 	Mux471;
output 	Mux44;
output 	Mux441;
output 	Mux46;
output 	Mux461;
output 	Mux42;
output 	Mux421;
output 	Mux43;
output 	Mux431;
output 	Mux35;
output 	Mux351;
output 	Mux37;
output 	Mux371;
output 	Mux55;
output 	Mux551;
output 	Mux56;
output 	Mux561;
output 	Mux41;
output 	Mux411;
output 	Mux38;
output 	Mux381;
output 	Mux29;
output 	Mux291;
output 	Mux27;
output 	Mux271;
output 	Mux28;
output 	Mux281;
output 	Mux23;
output 	Mux231;
output 	Mux24;
output 	Mux241;
output 	Mux25;
output 	Mux251;
output 	Mux26;
output 	Mux261;
output 	Mux15;
output 	Mux1510;
output 	Mux16;
output 	Mux165;
output 	Mux17;
output 	Mux171;
output 	Mux18;
output 	Mux181;
output 	Mux20;
output 	Mux201;
output 	Mux19;
output 	Mux191;
output 	Mux21;
output 	Mux211;
output 	Mux22;
output 	Mux221;
output 	Mux13;
output 	Mux131;
output 	Mux14;
output 	Mux1410;
output 	Mux11;
output 	Mux111;
output 	Mux12;
output 	Mux121;
output 	Mux9;
output 	Mux91;
output 	Mux10;
output 	Mux101;
output 	Mux7;
output 	Mux71;
output 	Mux8;
output 	Mux81;
output 	Mux0;
output 	Mux01;
output 	Mux1;
output 	Mux110;
output 	Mux2;
output 	Mux210;
output 	Mux5;
output 	Mux510;
output 	Mux6;
output 	Mux64;
output 	Mux3;
output 	Mux310;
output 	Mux4;
output 	Mux410;
input 	CLK;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Mux30~4_combout ;
wire \Mux30~14_combout ;
wire \reg_file[4][0]~q ;
wire \Mux63~12_combout ;
wire \Mux31~12_combout ;
wire \reg_file[16][2]~q ;
wire \reg_file[8][2]~q ;
wire \Mux59~4_combout ;
wire \reg_file[8][4]~q ;
wire \Mux32~4_combout ;
wire \Mux33~4_combout ;
wire \Mux33~14_combout ;
wire \Mux34~4_combout ;
wire \Mux58~2_combout ;
wire \Mux50~12_combout ;
wire \Mux52~12_combout ;
wire \Mux54~12_combout ;
wire \Mux36~2_combout ;
wire \reg_file[24][27]~q ;
wire \Mux40~4_combout ;
wire \reg_file[16][18]~q ;
wire \Mux45~4_combout ;
wire \Mux45~12_combout ;
wire \reg_file[2][18]~q ;
wire \reg_file[18][24]~q ;
wire \reg_file[20][24]~q ;
wire \Mux47~2_combout ;
wire \reg_file[26][19]~q ;
wire \reg_file[20][17]~q ;
wire \Mux46~4_combout ;
wire \Mux43~2_combout ;
wire \reg_file[8][20]~q ;
wire \reg_file[18][28]~q ;
wire \Mux35~2_combout ;
wire \Mux35~12_combout ;
wire \Mux37~2_combout ;
wire \reg_file[24][26]~q ;
wire \Mux37~4_combout ;
wire \Mux38~4_combout ;
wire \Mux38~14_combout ;
wire \Mux29~4_combout ;
wire \Mux29~12_combout ;
wire \Mux29~14_combout ;
wire \Mux27~2_combout ;
wire \Mux27~12_combout ;
wire \Mux28~14_combout ;
wire \Mux23~14_combout ;
wire \Mux25~2_combout ;
wire \Mux15~12_combout ;
wire \Mux17~14_combout ;
wire \Mux18~12_combout ;
wire \Mux19~2_combout ;
wire \Mux19~12_combout ;
wire \Mux19~14_combout ;
wire \Mux21~12_combout ;
wire \Mux22~2_combout ;
wire \Mux22~14_combout ;
wire \Mux13~4_combout ;
wire \Mux13~12_combout ;
wire \Mux14~12_combout ;
wire \Mux14~14_combout ;
wire \Mux11~12_combout ;
wire \Mux11~14_combout ;
wire \Mux12~2_combout ;
wire \Mux7~2_combout ;
wire \Mux7~4_combout ;
wire \Mux7~12_combout ;
wire \Mux7~14_combout ;
wire \Mux0~2_combout ;
wire \Mux1~2_combout ;
wire \Mux1~12_combout ;
wire \Mux2~2_combout ;
wire \Mux6~2_combout ;
wire \Mux3~2_combout ;
wire \Mux3~4_combout ;
wire \reg_file[24][27]~feeder_combout ;
wire \reg_file[2][18]~feeder_combout ;
wire \reg_file[26][19]~feeder_combout ;
wire \reg_file[20][17]~feeder_combout ;
wire \reg_file[18][28]~feeder_combout ;
wire \reg_file[24][26]~feeder_combout ;
wire \reg_file_nxt[31][1]~64_combout ;
wire \Decoder0~14_combout ;
wire \Decoder0~15_combout ;
wire \reg_file[21][1]~q ;
wire \Decoder0~19_combout ;
wire \reg_file[29][1]~q ;
wire \Decoder0~16_combout ;
wire \Decoder0~18_combout ;
wire \reg_file[17][1]~q ;
wire \Decoder0~17_combout ;
wire \reg_file[25][1]~q ;
wire \Mux62~0_combout ;
wire \Mux62~1_combout ;
wire \reg_file[30][1]~feeder_combout ;
wire \Decoder0~22_combout ;
wire \Decoder0~25_combout ;
wire \reg_file[30][1]~q ;
wire \Decoder0~20_combout ;
wire \Decoder0~24_combout ;
wire \reg_file[18][1]~q ;
wire \Decoder0~23_combout ;
wire \reg_file[22][1]~q ;
wire \Mux62~2_combout ;
wire \Decoder0~21_combout ;
wire \reg_file[26][1]~q ;
wire \Mux62~3_combout ;
wire \Decoder0~26_combout ;
wire \reg_file[24][1]~q ;
wire \Decoder0~27_combout ;
wire \reg_file[20][1]~q ;
wire \Decoder0~28_combout ;
wire \reg_file[16][1]~q ;
wire \Mux62~4_combout ;
wire \Mux62~5_combout ;
wire \Mux62~6_combout ;
wire \reg_file[23][1]~feeder_combout ;
wire \Decoder0~30_combout ;
wire \reg_file[23][1]~q ;
wire \Decoder0~33_combout ;
wire \reg_file[31][1]~q ;
wire \Decoder0~31_combout ;
wire \reg_file[27][1]~q ;
wire \Decoder0~32_combout ;
wire \reg_file[19][1]~q ;
wire \Mux62~7_combout ;
wire \Mux62~8_combout ;
wire \Decoder0~47_combout ;
wire \reg_file[1][1]~q ;
wire \reg_file[3][1]~feeder_combout ;
wire \Decoder0~46_combout ;
wire \reg_file[3][1]~q ;
wire \Mux62~14_combout ;
wire \Decoder0~48_combout ;
wire \reg_file[2][1]~q ;
wire \Mux62~15_combout ;
wire \Decoder0~34_combout ;
wire \reg_file[9][1]~q ;
wire \Decoder0~37_combout ;
wire \reg_file[11][1]~q ;
wire \Decoder0~35_combout ;
wire \reg_file[10][1]~q ;
wire \Mux62~12_combout ;
wire \Mux62~13_combout ;
wire \Mux62~16_combout ;
wire \Decoder0~39_combout ;
wire \reg_file[13][1]~q ;
wire \Decoder0~40_combout ;
wire \reg_file[12][1]~q ;
wire \Mux62~17_combout ;
wire \Decoder0~38_combout ;
wire \reg_file[14][1]~q ;
wire \Decoder0~41_combout ;
wire \reg_file[15][1]~q ;
wire \Mux62~18_combout ;
wire \reg_file[7][1]~feeder_combout ;
wire \Decoder0~45_combout ;
wire \reg_file[7][1]~q ;
wire \Decoder0~42_combout ;
wire \reg_file[6][1]~q ;
wire \Decoder0~44_combout ;
wire \reg_file[4][1]~q ;
wire \reg_file[5][1]~feeder_combout ;
wire \Decoder0~43_combout ;
wire \reg_file[5][1]~q ;
wire \Mux62~10_combout ;
wire \Mux62~11_combout ;
wire \Mux30~0_combout ;
wire \Mux30~1_combout ;
wire \Mux30~7_combout ;
wire \Mux30~8_combout ;
wire \Mux30~2_combout ;
wire \Mux30~3_combout ;
wire \Decoder0~29_combout ;
wire \reg_file[28][1]~q ;
wire \Mux30~5_combout ;
wire \Mux30~6_combout ;
wire \Mux30~15_combout ;
wire \Mux30~12_combout ;
wire \Mux30~13_combout ;
wire \Mux30~16_combout ;
wire \Decoder0~36_combout ;
wire \reg_file[8][1]~q ;
wire \Mux30~10_combout ;
wire \Mux30~11_combout ;
wire \Mux30~17_combout ;
wire \Mux30~18_combout ;
wire \reg_file_nxt[31][0]~65_combout ;
wire \reg_file[31][0]~q ;
wire \reg_file[19][0]~q ;
wire \reg_file[23][0]~q ;
wire \Mux63~7_combout ;
wire \reg_file[27][0]~q ;
wire \Mux63~8_combout ;
wire \reg_file[25][0]~feeder_combout ;
wire \reg_file[25][0]~q ;
wire \reg_file[29][0]~q ;
wire \reg_file[17][0]~q ;
wire \reg_file[21][0]~feeder_combout ;
wire \reg_file[21][0]~q ;
wire \Mux63~0_combout ;
wire \Mux63~1_combout ;
wire \reg_file[20][0]~q ;
wire \reg_file[28][0]~q ;
wire \reg_file[16][0]~q ;
wire \reg_file[24][0]~feeder_combout ;
wire \reg_file[24][0]~q ;
wire \Mux63~4_combout ;
wire \Mux63~5_combout ;
wire \reg_file[22][0]~q ;
wire \reg_file[18][0]~q ;
wire \reg_file[26][0]~feeder_combout ;
wire \reg_file[26][0]~q ;
wire \Mux63~2_combout ;
wire \Mux63~3_combout ;
wire \Mux63~6_combout ;
wire \reg_file[14][0]~q ;
wire \reg_file[13][0]~q ;
wire \reg_file[12][0]~q ;
wire \Mux63~17_combout ;
wire \reg_file[15][0]~q ;
wire \Mux63~18_combout ;
wire \reg_file[6][0]~feeder_combout ;
wire \reg_file[6][0]~q ;
wire \reg_file[7][0]~feeder_combout ;
wire \reg_file[7][0]~q ;
wire \Mux63~13_combout ;
wire \reg_file[2][0]~q ;
wire \reg_file[3][0]~q ;
wire \reg_file[1][0]~q ;
wire \Mux63~14_combout ;
wire \Mux63~15_combout ;
wire \Mux63~16_combout ;
wire \reg_file[11][0]~q ;
wire \reg_file[9][0]~q ;
wire \reg_file[10][0]~q ;
wire \reg_file[8][0]~q ;
wire \Mux63~10_combout ;
wire \Mux63~11_combout ;
wire \Mux31~7_combout ;
wire \Mux31~8_combout ;
wire \Mux31~4_combout ;
wire \Mux31~5_combout ;
wire \Mux31~2_combout ;
wire \reg_file[30][0]~q ;
wire \Mux31~3_combout ;
wire \Mux31~6_combout ;
wire \Mux31~0_combout ;
wire \Mux31~1_combout ;
wire \Mux31~13_combout ;
wire \Mux31~14_combout ;
wire \Mux31~15_combout ;
wire \Mux31~16_combout ;
wire \Mux31~17_combout ;
wire \Mux31~18_combout ;
wire \reg_file[5][0]~q ;
wire \Mux31~10_combout ;
wire \Mux31~11_combout ;
wire \reg_file_nxt[31][3]~66_combout ;
wire \reg_file[31][3]~q ;
wire \reg_file[23][3]~q ;
wire \reg_file[27][3]~q ;
wire \reg_file[19][3]~q ;
wire \Mux60~7_combout ;
wire \Mux60~8_combout ;
wire \reg_file[29][3]~feeder_combout ;
wire \reg_file[29][3]~q ;
wire \reg_file[21][3]~q ;
wire \reg_file[25][3]~feeder_combout ;
wire \reg_file[25][3]~q ;
wire \reg_file[17][3]~feeder_combout ;
wire \reg_file[17][3]~q ;
wire \Mux60~0_combout ;
wire \Mux60~1_combout ;
wire \reg_file[30][3]~feeder_combout ;
wire \reg_file[30][3]~q ;
wire \reg_file[18][3]~q ;
wire \reg_file[22][3]~feeder_combout ;
wire \reg_file[22][3]~q ;
wire \Mux60~2_combout ;
wire \Mux60~3_combout ;
wire \reg_file[28][3]~feeder_combout ;
wire \reg_file[28][3]~q ;
wire \reg_file[16][3]~q ;
wire \reg_file[20][3]~feeder_combout ;
wire \reg_file[20][3]~q ;
wire \Mux60~4_combout ;
wire \Mux60~5_combout ;
wire \Mux60~6_combout ;
wire \reg_file[14][3]~q ;
wire \reg_file[13][3]~q ;
wire \reg_file[12][3]~q ;
wire \Mux60~17_combout ;
wire \reg_file[15][3]~q ;
wire \Mux60~18_combout ;
wire \reg_file[2][3]~q ;
wire \reg_file[1][3]~q ;
wire \reg_file[3][3]~q ;
wire \Mux60~14_combout ;
wire \Mux60~15_combout ;
wire \reg_file[9][3]~q ;
wire \reg_file[11][3]~q ;
wire \reg_file[8][3]~q ;
wire \reg_file[10][3]~q ;
wire \Mux60~12_combout ;
wire \Mux60~13_combout ;
wire \Mux60~16_combout ;
wire \reg_file[6][3]~feeder_combout ;
wire \reg_file[6][3]~q ;
wire \reg_file[7][3]~q ;
wire \reg_file[5][3]~q ;
wire \reg_file[4][3]~q ;
wire \Mux60~10_combout ;
wire \Mux60~11_combout ;
wire \reg_file_nxt[31][2]~67_combout ;
wire \reg_file[22][2]~q ;
wire \reg_file[18][2]~feeder_combout ;
wire \reg_file[18][2]~q ;
wire \reg_file[26][2]~feeder_combout ;
wire \reg_file[26][2]~q ;
wire \Mux61~2_combout ;
wire \Mux61~3_combout ;
wire \reg_file[20][2]~q ;
wire \reg_file[24][2]~q ;
wire \Mux61~4_combout ;
wire \Mux61~5_combout ;
wire \Mux61~6_combout ;
wire \reg_file[23][2]~q ;
wire \reg_file[19][2]~q ;
wire \Mux61~7_combout ;
wire \reg_file[31][2]~feeder_combout ;
wire \reg_file[31][2]~q ;
wire \reg_file[27][2]~feeder_combout ;
wire \reg_file[27][2]~q ;
wire \Mux61~8_combout ;
wire \reg_file[25][2]~q ;
wire \reg_file[29][2]~feeder_combout ;
wire \reg_file[29][2]~q ;
wire \reg_file[17][2]~q ;
wire \reg_file[21][2]~feeder_combout ;
wire \reg_file[21][2]~q ;
wire \Mux61~0_combout ;
wire \Mux61~1_combout ;
wire \reg_file[10][2]~q ;
wire \Mux61~10_combout ;
wire \reg_file[9][2]~q ;
wire \reg_file[11][2]~q ;
wire \Mux61~11_combout ;
wire \reg_file[15][2]~q ;
wire \reg_file[14][2]~q ;
wire \reg_file[12][2]~q ;
wire \reg_file[13][2]~q ;
wire \Mux61~17_combout ;
wire \Mux61~18_combout ;
wire \reg_file[7][2]~q ;
wire \reg_file[4][2]~q ;
wire \reg_file[5][2]~q ;
wire \Mux61~12_combout ;
wire \Mux61~13_combout ;
wire \reg_file[2][2]~q ;
wire \reg_file[1][2]~q ;
wire \reg_file[3][2]~feeder_combout ;
wire \reg_file[3][2]~q ;
wire \Mux61~14_combout ;
wire \Mux61~15_combout ;
wire \Mux61~16_combout ;
wire \reg_file_nxt[31][4]~68_combout ;
wire \reg_file[27][4]~feeder_combout ;
wire \reg_file[27][4]~q ;
wire \reg_file[23][4]~q ;
wire \reg_file[19][4]~q ;
wire \Mux59~7_combout ;
wire \reg_file[31][4]~q ;
wire \Mux59~8_combout ;
wire \reg_file[22][4]~feeder_combout ;
wire \reg_file[22][4]~q ;
wire \reg_file[30][4]~q ;
wire \reg_file[26][4]~q ;
wire \reg_file[18][4]~q ;
wire \Mux59~2_combout ;
wire \Mux59~3_combout ;
wire \reg_file[28][4]~q ;
wire \reg_file[20][4]~q ;
wire \Mux59~5_combout ;
wire \Mux59~6_combout ;
wire \reg_file[29][4]~feeder_combout ;
wire \reg_file[29][4]~q ;
wire \reg_file[17][4]~q ;
wire \reg_file[21][4]~feeder_combout ;
wire \reg_file[21][4]~q ;
wire \Mux59~0_combout ;
wire \reg_file[25][4]~q ;
wire \Mux59~1_combout ;
wire \reg_file[10][4]~q ;
wire \Mux59~10_combout ;
wire \reg_file[9][4]~q ;
wire \reg_file[11][4]~q ;
wire \Mux59~11_combout ;
wire \reg_file[4][4]~q ;
wire \reg_file[5][4]~q ;
wire \Mux59~12_combout ;
wire \reg_file[7][4]~q ;
wire \Mux59~13_combout ;
wire \reg_file[2][4]~feeder_combout ;
wire \reg_file[2][4]~q ;
wire \reg_file[1][4]~q ;
wire \Mux59~14_combout ;
wire \Mux59~15_combout ;
wire \Mux59~16_combout ;
wire \reg_file[14][4]~q ;
wire \reg_file[12][4]~q ;
wire \reg_file[13][4]~q ;
wire \Mux59~17_combout ;
wire \reg_file[15][4]~q ;
wire \Mux59~18_combout ;
wire \reg_file_nxt[31][31]~69_combout ;
wire \reg_file[21][31]~q ;
wire \reg_file[29][31]~feeder_combout ;
wire \reg_file[29][31]~q ;
wire \reg_file[17][31]~q ;
wire \reg_file[25][31]~feeder_combout ;
wire \reg_file[25][31]~q ;
wire \Mux32~0_combout ;
wire \Mux32~1_combout ;
wire \reg_file[24][31]~q ;
wire \reg_file[28][31]~feeder_combout ;
wire \reg_file[28][31]~q ;
wire \Mux32~5_combout ;
wire \reg_file[18][31]~q ;
wire \Mux32~2_combout ;
wire \reg_file[30][31]~q ;
wire \reg_file[26][31]~q ;
wire \Mux32~3_combout ;
wire \Mux32~6_combout ;
wire \reg_file[23][31]~feeder_combout ;
wire \reg_file[23][31]~q ;
wire \reg_file[27][31]~q ;
wire \reg_file[19][31]~q ;
wire \Mux32~7_combout ;
wire \reg_file[31][31]~q ;
wire \Mux32~8_combout ;
wire \reg_file[14][31]~q ;
wire \reg_file[15][31]~q ;
wire \reg_file[12][31]~q ;
wire \reg_file[13][31]~q ;
wire \Mux32~17_combout ;
wire \Mux32~18_combout ;
wire \reg_file[7][31]~q ;
wire \reg_file[4][31]~q ;
wire \reg_file[5][31]~q ;
wire \Mux32~10_combout ;
wire \reg_file[6][31]~feeder_combout ;
wire \reg_file[6][31]~q ;
wire \Mux32~11_combout ;
wire \reg_file[2][31]~q ;
wire \reg_file[1][31]~q ;
wire \reg_file[3][31]~q ;
wire \Mux32~14_combout ;
wire \Mux32~15_combout ;
wire \reg_file[10][31]~q ;
wire \reg_file[8][31]~q ;
wire \Mux32~12_combout ;
wire \reg_file[11][31]~q ;
wire \reg_file[9][31]~q ;
wire \Mux32~13_combout ;
wire \Mux32~16_combout ;
wire \reg_file_nxt[31][30]~70_combout ;
wire \reg_file[31][30]~q ;
wire \reg_file[27][30]~q ;
wire \reg_file[23][30]~q ;
wire \reg_file[19][30]~q ;
wire \Mux33~7_combout ;
wire \Mux33~8_combout ;
wire \reg_file[25][30]~q ;
wire \reg_file[29][30]~q ;
wire \reg_file[17][30]~q ;
wire \reg_file[21][30]~feeder_combout ;
wire \reg_file[21][30]~q ;
wire \Mux33~0_combout ;
wire \Mux33~1_combout ;
wire \reg_file[18][30]~q ;
wire \reg_file[26][30]~q ;
wire \Mux33~2_combout ;
wire \reg_file[30][30]~q ;
wire \reg_file[22][30]~q ;
wire \Mux33~3_combout ;
wire \reg_file[28][30]~feeder_combout ;
wire \reg_file[28][30]~q ;
wire \reg_file[20][30]~q ;
wire \Mux33~5_combout ;
wire \Mux33~6_combout ;
wire \reg_file[6][30]~q ;
wire \reg_file[5][30]~q ;
wire \reg_file[4][30]~q ;
wire \Mux33~12_combout ;
wire \Mux33~13_combout ;
wire \reg_file[2][30]~q ;
wire \Mux33~15_combout ;
wire \Mux33~16_combout ;
wire \reg_file[14][30]~q ;
wire \reg_file[12][30]~q ;
wire \reg_file[13][30]~q ;
wire \Mux33~17_combout ;
wire \reg_file[15][30]~q ;
wire \Mux33~18_combout ;
wire \reg_file[11][30]~q ;
wire \reg_file[9][30]~q ;
wire \reg_file[8][30]~q ;
wire \reg_file[10][30]~q ;
wire \Mux33~10_combout ;
wire \Mux33~11_combout ;
wire \reg_file_nxt[31][29]~71_combout ;
wire \reg_file[27][29]~q ;
wire \reg_file[19][29]~q ;
wire \Mux34~7_combout ;
wire \reg_file[23][29]~q ;
wire \reg_file[31][29]~q ;
wire \Mux34~8_combout ;
wire \reg_file[29][29]~feeder_combout ;
wire \reg_file[29][29]~q ;
wire \reg_file[17][29]~q ;
wire \reg_file[25][29]~feeder_combout ;
wire \reg_file[25][29]~q ;
wire \Mux34~0_combout ;
wire \reg_file[21][29]~q ;
wire \Mux34~1_combout ;
wire \reg_file[26][29]~q ;
wire \reg_file[30][29]~q ;
wire \reg_file[18][29]~q ;
wire \reg_file[22][29]~q ;
wire \Mux34~2_combout ;
wire \Mux34~3_combout ;
wire \reg_file[28][29]~q ;
wire \reg_file[24][29]~q ;
wire \Mux34~5_combout ;
wire \Mux34~6_combout ;
wire \reg_file[14][29]~feeder_combout ;
wire \reg_file[14][29]~q ;
wire \reg_file[12][29]~q ;
wire \reg_file[13][29]~q ;
wire \Mux34~17_combout ;
wire \reg_file[15][29]~feeder_combout ;
wire \reg_file[15][29]~q ;
wire \Mux34~18_combout ;
wire \reg_file[2][29]~q ;
wire \reg_file[1][29]~q ;
wire \reg_file[3][29]~q ;
wire \Mux34~14_combout ;
wire \Mux34~15_combout ;
wire \reg_file[11][29]~q ;
wire \reg_file[10][29]~q ;
wire \reg_file[8][29]~q ;
wire \Mux34~12_combout ;
wire \Mux34~13_combout ;
wire \Mux34~16_combout ;
wire \reg_file[4][29]~q ;
wire \reg_file[5][29]~q ;
wire \Mux34~10_combout ;
wire \reg_file[6][29]~q ;
wire \reg_file[7][29]~q ;
wire \Mux34~11_combout ;
wire \reg_file_nxt[31][5]~72_combout ;
wire \reg_file[30][5]~q ;
wire \reg_file[26][5]~q ;
wire \Mux58~3_combout ;
wire \reg_file[24][5]~q ;
wire \reg_file[20][5]~q ;
wire \reg_file[16][5]~q ;
wire \Mux58~4_combout ;
wire \Mux58~5_combout ;
wire \Mux58~6_combout ;
wire \reg_file[25][5]~q ;
wire \reg_file[17][5]~q ;
wire \Mux58~0_combout ;
wire \reg_file[21][5]~feeder_combout ;
wire \reg_file[21][5]~q ;
wire \reg_file[29][5]~feeder_combout ;
wire \reg_file[29][5]~q ;
wire \Mux58~1_combout ;
wire \reg_file[23][5]~feeder_combout ;
wire \reg_file[23][5]~q ;
wire \reg_file[31][5]~feeder_combout ;
wire \reg_file[31][5]~q ;
wire \reg_file[27][5]~q ;
wire \reg_file[19][5]~q ;
wire \Mux58~7_combout ;
wire \Mux58~8_combout ;
wire \reg_file[6][5]~feeder_combout ;
wire \reg_file[6][5]~q ;
wire \reg_file[7][5]~q ;
wire \reg_file[4][5]~q ;
wire \reg_file[5][5]~q ;
wire \Mux58~10_combout ;
wire \Mux58~11_combout ;
wire \reg_file[1][5]~q ;
wire \reg_file[3][5]~q ;
wire \Mux58~14_combout ;
wire \Mux58~15_combout ;
wire \reg_file[9][5]~feeder_combout ;
wire \reg_file[9][5]~q ;
wire \reg_file[11][5]~q ;
wire \reg_file[10][5]~q ;
wire \reg_file[8][5]~q ;
wire \Mux58~12_combout ;
wire \Mux58~13_combout ;
wire \Mux58~16_combout ;
wire \reg_file[13][5]~q ;
wire \reg_file[12][5]~q ;
wire \Mux58~17_combout ;
wire \reg_file[14][5]~feeder_combout ;
wire \reg_file[14][5]~q ;
wire \reg_file[15][5]~q ;
wire \Mux58~18_combout ;
wire \reg_file_nxt[31][15]~73_combout ;
wire \reg_file[29][15]~feeder_combout ;
wire \reg_file[29][15]~q ;
wire \reg_file[21][15]~q ;
wire \reg_file[17][15]~q ;
wire \reg_file[25][15]~q ;
wire \Mux48~0_combout ;
wire \Mux48~1_combout ;
wire \reg_file[27][15]~q ;
wire \reg_file[19][15]~q ;
wire \Mux48~7_combout ;
wire \reg_file[31][15]~q ;
wire \reg_file[23][15]~feeder_combout ;
wire \reg_file[23][15]~q ;
wire \Mux48~8_combout ;
wire \reg_file[28][15]~q ;
wire \reg_file[24][15]~q ;
wire \reg_file[20][15]~q ;
wire \reg_file[16][15]~q ;
wire \Mux48~4_combout ;
wire \Mux48~5_combout ;
wire \reg_file[22][15]~q ;
wire \reg_file[18][15]~q ;
wire \Mux48~2_combout ;
wire \reg_file[30][15]~q ;
wire \reg_file[26][15]~q ;
wire \Mux48~3_combout ;
wire \Mux48~6_combout ;
wire \reg_file[2][15]~feeder_combout ;
wire \reg_file[2][15]~q ;
wire \reg_file[3][15]~feeder_combout ;
wire \reg_file[3][15]~q ;
wire \reg_file[1][15]~q ;
wire \Mux48~14_combout ;
wire \Mux48~15_combout ;
wire \reg_file[9][15]~q ;
wire \reg_file[11][15]~q ;
wire \reg_file[10][15]~q ;
wire \reg_file[8][15]~q ;
wire \Mux48~12_combout ;
wire \Mux48~13_combout ;
wire \Mux48~16_combout ;
wire \reg_file[6][15]~feeder_combout ;
wire \reg_file[6][15]~q ;
wire \reg_file[5][15]~q ;
wire \reg_file[4][15]~q ;
wire \Mux48~10_combout ;
wire \reg_file[7][15]~q ;
wire \Mux48~11_combout ;
wire \reg_file[12][15]~q ;
wire \reg_file[13][15]~q ;
wire \Mux48~17_combout ;
wire \reg_file[14][15]~q ;
wire \reg_file[15][15]~q ;
wire \Mux48~18_combout ;
wire \reg_file_nxt[31][14]~74_combout ;
wire \reg_file[18][14]~q ;
wire \reg_file[26][14]~feeder_combout ;
wire \reg_file[26][14]~q ;
wire \Mux49~2_combout ;
wire \reg_file[22][14]~q ;
wire \Mux49~3_combout ;
wire \reg_file[28][14]~q ;
wire \reg_file[20][14]~q ;
wire \reg_file[16][14]~q ;
wire \reg_file[24][14]~q ;
wire \Mux49~4_combout ;
wire \Mux49~5_combout ;
wire \Mux49~6_combout ;
wire \reg_file[23][14]~q ;
wire \reg_file[19][14]~q ;
wire \Mux49~7_combout ;
wire \reg_file[27][14]~feeder_combout ;
wire \reg_file[27][14]~q ;
wire \reg_file[31][14]~feeder_combout ;
wire \reg_file[31][14]~q ;
wire \Mux49~8_combout ;
wire \reg_file[25][14]~feeder_combout ;
wire \reg_file[25][14]~q ;
wire \reg_file[29][14]~q ;
wire \reg_file[17][14]~q ;
wire \reg_file[21][14]~q ;
wire \Mux49~0_combout ;
wire \Mux49~1_combout ;
wire \reg_file[13][14]~q ;
wire \reg_file[12][14]~q ;
wire \Mux49~17_combout ;
wire \reg_file[15][14]~q ;
wire \reg_file[14][14]~feeder_combout ;
wire \reg_file[14][14]~q ;
wire \Mux49~18_combout ;
wire \reg_file[10][14]~q ;
wire \Mux49~10_combout ;
wire \reg_file[9][14]~feeder_combout ;
wire \reg_file[9][14]~q ;
wire \reg_file[11][14]~q ;
wire \Mux49~11_combout ;
wire \reg_file[6][14]~feeder_combout ;
wire \reg_file[6][14]~q ;
wire \reg_file[7][14]~q ;
wire \reg_file[4][14]~q ;
wire \reg_file[5][14]~q ;
wire \Mux49~12_combout ;
wire \Mux49~13_combout ;
wire \reg_file[2][14]~q ;
wire \reg_file[1][14]~q ;
wire \reg_file[3][14]~q ;
wire \Mux49~14_combout ;
wire \Mux49~15_combout ;
wire \Mux49~16_combout ;
wire \reg_file_nxt[31][13]~75_combout ;
wire \reg_file[30][13]~q ;
wire \reg_file[22][13]~feeder_combout ;
wire \reg_file[22][13]~q ;
wire \reg_file[18][13]~q ;
wire \Mux50~2_combout ;
wire \Mux50~3_combout ;
wire \reg_file[24][13]~q ;
wire \reg_file[20][13]~q ;
wire \Mux50~4_combout ;
wire \Mux50~5_combout ;
wire \Mux50~6_combout ;
wire \reg_file[25][13]~q ;
wire \Mux50~0_combout ;
wire \reg_file[21][13]~q ;
wire \reg_file[29][13]~feeder_combout ;
wire \reg_file[29][13]~q ;
wire \Mux50~1_combout ;
wire \reg_file[31][13]~q ;
wire \reg_file[23][13]~q ;
wire \reg_file[27][13]~q ;
wire \reg_file[19][13]~q ;
wire \Mux50~7_combout ;
wire \Mux50~8_combout ;
wire \reg_file[6][13]~feeder_combout ;
wire \reg_file[6][13]~q ;
wire \reg_file[7][13]~q ;
wire \reg_file[5][13]~feeder_combout ;
wire \reg_file[5][13]~q ;
wire \reg_file[4][13]~q ;
wire \Mux50~10_combout ;
wire \Mux50~11_combout ;
wire \reg_file[13][13]~q ;
wire \Mux50~17_combout ;
wire \reg_file[15][13]~q ;
wire \reg_file[14][13]~q ;
wire \Mux50~18_combout ;
wire \reg_file[2][13]~q ;
wire \reg_file[3][13]~q ;
wire \reg_file[1][13]~q ;
wire \Mux50~14_combout ;
wire \Mux50~15_combout ;
wire \reg_file[11][13]~q ;
wire \reg_file[9][13]~q ;
wire \Mux50~13_combout ;
wire \Mux50~16_combout ;
wire \reg_file_nxt[31][12]~76_combout ;
wire \reg_file[27][12]~feeder_combout ;
wire \reg_file[27][12]~q ;
wire \reg_file[19][12]~q ;
wire \reg_file[23][12]~q ;
wire \Mux51~7_combout ;
wire \reg_file[31][12]~feeder_combout ;
wire \reg_file[31][12]~q ;
wire \Mux51~8_combout ;
wire \reg_file[30][12]~q ;
wire \reg_file[22][12]~feeder_combout ;
wire \reg_file[22][12]~q ;
wire \reg_file[18][12]~q ;
wire \reg_file[26][12]~feeder_combout ;
wire \reg_file[26][12]~q ;
wire \Mux51~2_combout ;
wire \Mux51~3_combout ;
wire \reg_file[28][12]~feeder_combout ;
wire \reg_file[28][12]~q ;
wire \reg_file[20][12]~q ;
wire \reg_file[16][12]~q ;
wire \reg_file[24][12]~q ;
wire \Mux51~4_combout ;
wire \Mux51~5_combout ;
wire \Mux51~6_combout ;
wire \reg_file[29][12]~feeder_combout ;
wire \reg_file[29][12]~q ;
wire \reg_file[25][12]~feeder_combout ;
wire \reg_file[25][12]~q ;
wire \reg_file[21][12]~feeder_combout ;
wire \reg_file[21][12]~q ;
wire \reg_file[17][12]~q ;
wire \Mux51~0_combout ;
wire \Mux51~1_combout ;
wire \reg_file[11][12]~q ;
wire \reg_file[8][12]~q ;
wire \reg_file[10][12]~q ;
wire \Mux51~10_combout ;
wire \reg_file[9][12]~q ;
wire \Mux51~11_combout ;
wire \reg_file[3][12]~q ;
wire \reg_file[1][12]~q ;
wire \Mux51~14_combout ;
wire \reg_file[2][12]~feeder_combout ;
wire \reg_file[2][12]~q ;
wire \Mux51~15_combout ;
wire \reg_file[4][12]~q ;
wire \reg_file[5][12]~q ;
wire \Mux51~12_combout ;
wire \reg_file[7][12]~feeder_combout ;
wire \reg_file[7][12]~q ;
wire \Mux51~13_combout ;
wire \Mux51~16_combout ;
wire \reg_file[12][12]~q ;
wire \reg_file[13][12]~q ;
wire \Mux51~17_combout ;
wire \reg_file[14][12]~feeder_combout ;
wire \reg_file[14][12]~q ;
wire \reg_file[15][12]~q ;
wire \Mux51~18_combout ;
wire \reg_file_nxt[31][11]~77_combout ;
wire \reg_file[23][11]~feeder_combout ;
wire \reg_file[23][11]~q ;
wire \reg_file[31][11]~q ;
wire \reg_file[27][11]~q ;
wire \reg_file[19][11]~q ;
wire \Mux52~7_combout ;
wire \Mux52~8_combout ;
wire \reg_file[25][11]~q ;
wire \Mux52~0_combout ;
wire \reg_file[21][11]~q ;
wire \reg_file[29][11]~q ;
wire \Mux52~1_combout ;
wire \reg_file[28][11]~q ;
wire \reg_file[24][11]~q ;
wire \reg_file[16][11]~q ;
wire \reg_file[20][11]~q ;
wire \Mux52~4_combout ;
wire \Mux52~5_combout ;
wire \reg_file[26][11]~q ;
wire \reg_file[30][11]~q ;
wire \reg_file[18][11]~q ;
wire \reg_file[22][11]~feeder_combout ;
wire \reg_file[22][11]~q ;
wire \Mux52~2_combout ;
wire \Mux52~3_combout ;
wire \Mux52~6_combout ;
wire \reg_file[11][11]~q ;
wire \reg_file[9][11]~q ;
wire \Mux52~13_combout ;
wire \reg_file[2][11]~q ;
wire \reg_file[3][11]~q ;
wire \reg_file[1][11]~q ;
wire \Mux52~14_combout ;
wire \Mux52~15_combout ;
wire \Mux52~16_combout ;
wire \reg_file[6][11]~feeder_combout ;
wire \reg_file[6][11]~q ;
wire \reg_file[4][11]~q ;
wire \reg_file[5][11]~q ;
wire \Mux52~10_combout ;
wire \reg_file[7][11]~q ;
wire \Mux52~11_combout ;
wire \reg_file[13][11]~q ;
wire \reg_file[12][11]~q ;
wire \Mux52~17_combout ;
wire \reg_file[14][11]~q ;
wire \reg_file[15][11]~q ;
wire \Mux52~18_combout ;
wire \reg_file_nxt[31][10]~78_combout ;
wire \reg_file[29][10]~q ;
wire \reg_file[25][10]~q ;
wire \reg_file[17][10]~q ;
wire \reg_file[21][10]~feeder_combout ;
wire \reg_file[21][10]~q ;
wire \Mux53~0_combout ;
wire \Mux53~1_combout ;
wire \reg_file[18][10]~q ;
wire \reg_file[26][10]~q ;
wire \Mux53~2_combout ;
wire \reg_file[30][10]~q ;
wire \reg_file[22][10]~q ;
wire \Mux53~3_combout ;
wire \reg_file[24][10]~q ;
wire \reg_file[16][10]~q ;
wire \Mux53~4_combout ;
wire \reg_file[20][10]~q ;
wire \Mux53~5_combout ;
wire \Mux53~6_combout ;
wire \reg_file[27][10]~feeder_combout ;
wire \reg_file[27][10]~q ;
wire \reg_file[31][10]~q ;
wire \reg_file[23][10]~q ;
wire \reg_file[19][10]~q ;
wire \Mux53~7_combout ;
wire \Mux53~8_combout ;
wire \reg_file[12][10]~q ;
wire \reg_file[13][10]~q ;
wire \Mux53~17_combout ;
wire \reg_file[15][10]~q ;
wire \reg_file[14][10]~feeder_combout ;
wire \reg_file[14][10]~q ;
wire \Mux53~18_combout ;
wire \reg_file[8][10]~q ;
wire \reg_file[10][10]~q ;
wire \Mux53~10_combout ;
wire \reg_file[9][10]~q ;
wire \reg_file[11][10]~q ;
wire \Mux53~11_combout ;
wire \reg_file[2][10]~q ;
wire \reg_file[1][10]~q ;
wire \reg_file[3][10]~q ;
wire \Mux53~14_combout ;
wire \Mux53~15_combout ;
wire \reg_file[6][10]~q ;
wire \reg_file[7][10]~q ;
wire \reg_file[5][10]~q ;
wire \reg_file[4][10]~q ;
wire \Mux53~12_combout ;
wire \Mux53~13_combout ;
wire \Mux53~16_combout ;
wire \reg_file_nxt[31][9]~79_combout ;
wire \reg_file[24][9]~q ;
wire \reg_file[16][9]~feeder_combout ;
wire \reg_file[16][9]~q ;
wire \reg_file[20][9]~feeder_combout ;
wire \reg_file[20][9]~q ;
wire \Mux54~4_combout ;
wire \reg_file[28][9]~q ;
wire \Mux54~5_combout ;
wire \reg_file[26][9]~q ;
wire \reg_file[30][9]~feeder_combout ;
wire \reg_file[30][9]~q ;
wire \reg_file[18][9]~q ;
wire \reg_file[22][9]~q ;
wire \Mux54~2_combout ;
wire \Mux54~3_combout ;
wire \Mux54~6_combout ;
wire \reg_file[29][9]~q ;
wire \reg_file[21][9]~q ;
wire \reg_file[17][9]~q ;
wire \reg_file[25][9]~q ;
wire \Mux54~0_combout ;
wire \Mux54~1_combout ;
wire \reg_file[27][9]~q ;
wire \Mux54~7_combout ;
wire \reg_file[23][9]~q ;
wire \reg_file[31][9]~q ;
wire \Mux54~8_combout ;
wire \reg_file[12][9]~q ;
wire \reg_file[13][9]~q ;
wire \Mux54~17_combout ;
wire \reg_file[14][9]~q ;
wire \reg_file[15][9]~q ;
wire \Mux54~18_combout ;
wire \reg_file[2][9]~feeder_combout ;
wire \reg_file[2][9]~q ;
wire \reg_file[1][9]~q ;
wire \reg_file[3][9]~q ;
wire \Mux54~14_combout ;
wire \Mux54~15_combout ;
wire \reg_file[11][9]~feeder_combout ;
wire \reg_file[11][9]~q ;
wire \reg_file[9][9]~q ;
wire \Mux54~13_combout ;
wire \Mux54~16_combout ;
wire \reg_file[6][9]~feeder_combout ;
wire \reg_file[6][9]~q ;
wire \reg_file[5][9]~q ;
wire \reg_file[4][9]~q ;
wire \Mux54~10_combout ;
wire \reg_file[7][9]~q ;
wire \Mux54~11_combout ;
wire \reg_file_nxt[31][6]~80_combout ;
wire \reg_file[25][6]~q ;
wire \reg_file[17][6]~q ;
wire \Mux57~0_combout ;
wire \reg_file[29][6]~feeder_combout ;
wire \reg_file[29][6]~q ;
wire \Mux57~1_combout ;
wire \reg_file[23][6]~q ;
wire \reg_file[19][6]~q ;
wire \Mux57~7_combout ;
wire \reg_file[31][6]~q ;
wire \reg_file[27][6]~feeder_combout ;
wire \reg_file[27][6]~q ;
wire \Mux57~8_combout ;
wire \reg_file[22][6]~q ;
wire \reg_file[18][6]~q ;
wire \reg_file[26][6]~feeder_combout ;
wire \reg_file[26][6]~q ;
wire \Mux57~2_combout ;
wire \Mux57~3_combout ;
wire \reg_file[28][6]~q ;
wire \reg_file[16][6]~q ;
wire \reg_file[24][6]~feeder_combout ;
wire \reg_file[24][6]~q ;
wire \Mux57~4_combout ;
wire \Mux57~5_combout ;
wire \Mux57~6_combout ;
wire \reg_file[1][6]~q ;
wire \reg_file[3][6]~feeder_combout ;
wire \reg_file[3][6]~q ;
wire \Mux57~14_combout ;
wire \reg_file[2][6]~q ;
wire \Mux57~15_combout ;
wire \reg_file[6][6]~q ;
wire \reg_file[7][6]~q ;
wire \reg_file[5][6]~q ;
wire \reg_file[4][6]~q ;
wire \Mux57~12_combout ;
wire \Mux57~13_combout ;
wire \Mux57~16_combout ;
wire \reg_file[9][6]~q ;
wire \reg_file[11][6]~q ;
wire \reg_file[10][6]~q ;
wire \reg_file[8][6]~q ;
wire \Mux57~10_combout ;
wire \Mux57~11_combout ;
wire \reg_file[15][6]~q ;
wire \reg_file[14][6]~feeder_combout ;
wire \reg_file[14][6]~q ;
wire \reg_file[13][6]~q ;
wire \reg_file[12][6]~q ;
wire \Mux57~17_combout ;
wire \Mux57~18_combout ;
wire \reg_file_nxt[31][27]~81_combout ;
wire \reg_file[26][27]~q ;
wire \reg_file[30][27]~q ;
wire \Mux36~3_combout ;
wire \reg_file[28][27]~q ;
wire \reg_file[20][27]~q ;
wire \Mux36~4_combout ;
wire \Mux36~5_combout ;
wire \Mux36~6_combout ;
wire \reg_file[29][27]~feeder_combout ;
wire \reg_file[29][27]~q ;
wire \reg_file[21][27]~q ;
wire \reg_file[17][27]~q ;
wire \Mux36~0_combout ;
wire \Mux36~1_combout ;
wire \reg_file[27][27]~q ;
wire \reg_file[19][27]~q ;
wire \Mux36~7_combout ;
wire \reg_file[23][27]~feeder_combout ;
wire \reg_file[23][27]~q ;
wire \reg_file[31][27]~feeder_combout ;
wire \reg_file[31][27]~q ;
wire \Mux36~8_combout ;
wire \reg_file[15][27]~q ;
wire \reg_file[13][27]~q ;
wire \reg_file[12][27]~q ;
wire \Mux36~17_combout ;
wire \reg_file[14][27]~feeder_combout ;
wire \reg_file[14][27]~q ;
wire \Mux36~18_combout ;
wire \reg_file[1][27]~q ;
wire \reg_file[3][27]~feeder_combout ;
wire \reg_file[3][27]~q ;
wire \Mux36~14_combout ;
wire \reg_file[2][27]~feeder_combout ;
wire \reg_file[2][27]~q ;
wire \Mux36~15_combout ;
wire \reg_file[9][27]~q ;
wire \reg_file[11][27]~q ;
wire \reg_file[8][27]~q ;
wire \reg_file[10][27]~q ;
wire \Mux36~12_combout ;
wire \Mux36~13_combout ;
wire \Mux36~16_combout ;
wire \reg_file[7][27]~q ;
wire \reg_file[6][27]~q ;
wire \reg_file[5][27]~q ;
wire \reg_file[4][27]~q ;
wire \Mux36~10_combout ;
wire \Mux36~11_combout ;
wire \reg_file_nxt[31][23]~82_combout ;
wire \reg_file[21][23]~feeder_combout ;
wire \reg_file[21][23]~q ;
wire \reg_file[25][23]~q ;
wire \Mux40~0_combout ;
wire \reg_file[29][23]~feeder_combout ;
wire \reg_file[29][23]~q ;
wire \Mux40~1_combout ;
wire \reg_file[18][23]~q ;
wire \reg_file[22][23]~q ;
wire \Mux40~2_combout ;
wire \reg_file[30][23]~q ;
wire \reg_file[26][23]~feeder_combout ;
wire \reg_file[26][23]~q ;
wire \Mux40~3_combout ;
wire \reg_file[28][23]~q ;
wire \reg_file[24][23]~q ;
wire \Mux40~5_combout ;
wire \Mux40~6_combout ;
wire \reg_file[27][23]~q ;
wire \reg_file[19][23]~q ;
wire \Mux40~7_combout ;
wire \reg_file[23][23]~q ;
wire \reg_file[31][23]~feeder_combout ;
wire \reg_file[31][23]~q ;
wire \Mux40~8_combout ;
wire \reg_file[14][23]~q ;
wire \reg_file[15][23]~q ;
wire \reg_file[12][23]~q ;
wire \reg_file[13][23]~q ;
wire \Mux40~17_combout ;
wire \Mux40~18_combout ;
wire \reg_file[6][23]~feeder_combout ;
wire \reg_file[6][23]~q ;
wire \reg_file[7][23]~feeder_combout ;
wire \reg_file[7][23]~q ;
wire \reg_file[5][23]~q ;
wire \reg_file[4][23]~q ;
wire \Mux40~10_combout ;
wire \Mux40~11_combout ;
wire \reg_file[8][23]~q ;
wire \reg_file[10][23]~q ;
wire \Mux40~12_combout ;
wire \reg_file[11][23]~q ;
wire \Mux40~13_combout ;
wire \reg_file[2][23]~feeder_combout ;
wire \reg_file[2][23]~q ;
wire \reg_file[3][23]~q ;
wire \reg_file[1][23]~q ;
wire \Mux40~14_combout ;
wire \Mux40~15_combout ;
wire \Mux40~16_combout ;
wire \reg_file_nxt[31][18]~83_combout ;
wire \reg_file[30][18]~feeder_combout ;
wire \reg_file[30][18]~q ;
wire \reg_file[22][18]~feeder_combout ;
wire \reg_file[22][18]~q ;
wire \reg_file[18][18]~q ;
wire \reg_file[26][18]~q ;
wire \Mux45~2_combout ;
wire \Mux45~3_combout ;
wire \reg_file[20][18]~q ;
wire \reg_file[28][18]~q ;
wire \Mux45~5_combout ;
wire \Mux45~6_combout ;
wire \reg_file[23][18]~q ;
wire \reg_file[19][18]~q ;
wire \Mux45~7_combout ;
wire \reg_file[27][18]~q ;
wire \reg_file[31][18]~q ;
wire \Mux45~8_combout ;
wire \reg_file[25][18]~q ;
wire \reg_file[29][18]~feeder_combout ;
wire \reg_file[29][18]~q ;
wire \reg_file[17][18]~q ;
wire \reg_file[21][18]~feeder_combout ;
wire \reg_file[21][18]~q ;
wire \Mux45~0_combout ;
wire \Mux45~1_combout ;
wire \reg_file[7][18]~q ;
wire \reg_file[6][18]~q ;
wire \Mux45~13_combout ;
wire \reg_file[1][18]~q ;
wire \Mux45~14_combout ;
wire \Mux45~15_combout ;
wire \Mux45~16_combout ;
wire \reg_file[14][18]~feeder_combout ;
wire \reg_file[14][18]~q ;
wire \reg_file[15][18]~q ;
wire \reg_file[13][18]~q ;
wire \Mux45~17_combout ;
wire \Mux45~18_combout ;
wire \reg_file[11][18]~feeder_combout ;
wire \reg_file[11][18]~q ;
wire \reg_file[9][18]~q ;
wire \reg_file[8][18]~q ;
wire \reg_file[10][18]~q ;
wire \Mux45~10_combout ;
wire \Mux45~11_combout ;
wire \reg_file_nxt[31][24]~84_combout ;
wire \reg_file[29][24]~feeder_combout ;
wire \reg_file[29][24]~q ;
wire \reg_file[25][24]~q ;
wire \reg_file[17][24]~q ;
wire \reg_file[21][24]~feeder_combout ;
wire \reg_file[21][24]~q ;
wire \Mux39~0_combout ;
wire \Mux39~1_combout ;
wire \reg_file[28][24]~q ;
wire \reg_file[16][24]~q ;
wire \Mux39~4_combout ;
wire \Mux39~5_combout ;
wire \reg_file[26][24]~q ;
wire \Mux39~2_combout ;
wire \reg_file[22][24]~q ;
wire \Mux39~3_combout ;
wire \Mux39~6_combout ;
wire \reg_file[31][24]~feeder_combout ;
wire \reg_file[31][24]~q ;
wire \reg_file[27][24]~q ;
wire \reg_file[23][24]~q ;
wire \reg_file[19][24]~q ;
wire \Mux39~7_combout ;
wire \Mux39~8_combout ;
wire \reg_file[6][24]~q ;
wire \reg_file[7][24]~q ;
wire \reg_file[4][24]~q ;
wire \reg_file[5][24]~q ;
wire \Mux39~12_combout ;
wire \Mux39~13_combout ;
wire \reg_file[1][24]~q ;
wire \reg_file[3][24]~feeder_combout ;
wire \reg_file[3][24]~q ;
wire \Mux39~14_combout ;
wire \reg_file[2][24]~q ;
wire \Mux39~15_combout ;
wire \Mux39~16_combout ;
wire \reg_file[11][24]~q ;
wire \reg_file[9][24]~q ;
wire \reg_file[8][24]~q ;
wire \reg_file[10][24]~q ;
wire \Mux39~10_combout ;
wire \Mux39~11_combout ;
wire \reg_file[15][24]~q ;
wire \reg_file[14][24]~feeder_combout ;
wire \reg_file[14][24]~q ;
wire \reg_file[12][24]~q ;
wire \reg_file[13][24]~q ;
wire \Mux39~17_combout ;
wire \Mux39~18_combout ;
wire \reg_file_nxt[31][16]~85_combout ;
wire \reg_file[25][16]~q ;
wire \reg_file[29][16]~feeder_combout ;
wire \reg_file[29][16]~q ;
wire \reg_file[17][16]~q ;
wire \Mux47~0_combout ;
wire \Mux47~1_combout ;
wire \reg_file[31][16]~feeder_combout ;
wire \reg_file[31][16]~q ;
wire \reg_file[27][16]~feeder_combout ;
wire \reg_file[27][16]~q ;
wire \reg_file[23][16]~q ;
wire \Mux47~7_combout ;
wire \Mux47~8_combout ;
wire \reg_file[28][16]~q ;
wire \reg_file[20][16]~q ;
wire \reg_file[24][16]~feeder_combout ;
wire \reg_file[24][16]~q ;
wire \reg_file[16][16]~q ;
wire \Mux47~4_combout ;
wire \Mux47~5_combout ;
wire \reg_file[30][16]~q ;
wire \reg_file[22][16]~feeder_combout ;
wire \reg_file[22][16]~q ;
wire \Mux47~3_combout ;
wire \Mux47~6_combout ;
wire \reg_file[1][16]~q ;
wire \Mux47~14_combout ;
wire \reg_file[2][16]~q ;
wire \Mux47~15_combout ;
wire \reg_file[6][16]~q ;
wire \reg_file[7][16]~q ;
wire \reg_file[4][16]~q ;
wire \reg_file[5][16]~q ;
wire \Mux47~12_combout ;
wire \Mux47~13_combout ;
wire \Mux47~16_combout ;
wire \reg_file[12][16]~q ;
wire \reg_file[13][16]~q ;
wire \Mux47~17_combout ;
wire \reg_file[14][16]~q ;
wire \reg_file[15][16]~feeder_combout ;
wire \reg_file[15][16]~q ;
wire \Mux47~18_combout ;
wire \reg_file[9][16]~feeder_combout ;
wire \reg_file[9][16]~q ;
wire \reg_file[8][16]~q ;
wire \reg_file[10][16]~q ;
wire \Mux47~10_combout ;
wire \reg_file[11][16]~feeder_combout ;
wire \reg_file[11][16]~q ;
wire \Mux47~11_combout ;
wire \reg_file_nxt[31][19]~86_combout ;
wire \reg_file[29][19]~feeder_combout ;
wire \reg_file[29][19]~q ;
wire \reg_file[21][19]~feeder_combout ;
wire \reg_file[21][19]~q ;
wire \reg_file[17][19]~q ;
wire \reg_file[25][19]~q ;
wire \Mux44~0_combout ;
wire \Mux44~1_combout ;
wire \reg_file[20][19]~feeder_combout ;
wire \reg_file[20][19]~q ;
wire \reg_file[16][19]~q ;
wire \Mux44~4_combout ;
wire \reg_file[28][19]~q ;
wire \Mux44~5_combout ;
wire \reg_file[22][19]~q ;
wire \reg_file[18][19]~q ;
wire \Mux44~2_combout ;
wire \reg_file[30][19]~q ;
wire \Mux44~3_combout ;
wire \Mux44~6_combout ;
wire \reg_file[19][19]~q ;
wire \reg_file[27][19]~q ;
wire \Mux44~7_combout ;
wire \reg_file[23][19]~feeder_combout ;
wire \reg_file[23][19]~q ;
wire \reg_file[31][19]~feeder_combout ;
wire \reg_file[31][19]~q ;
wire \Mux44~8_combout ;
wire \reg_file[6][19]~feeder_combout ;
wire \reg_file[6][19]~q ;
wire \reg_file[7][19]~q ;
wire \reg_file[4][19]~q ;
wire \reg_file[5][19]~q ;
wire \Mux44~10_combout ;
wire \Mux44~11_combout ;
wire \reg_file[15][19]~q ;
wire \reg_file[12][19]~q ;
wire \reg_file[13][19]~q ;
wire \Mux44~17_combout ;
wire \reg_file[14][19]~q ;
wire \Mux44~18_combout ;
wire \reg_file[3][19]~q ;
wire \reg_file[1][19]~q ;
wire \Mux44~14_combout ;
wire \reg_file[2][19]~feeder_combout ;
wire \reg_file[2][19]~q ;
wire \Mux44~15_combout ;
wire \reg_file[10][19]~q ;
wire \reg_file[8][19]~q ;
wire \Mux44~12_combout ;
wire \reg_file[9][19]~q ;
wire \Mux44~13_combout ;
wire \Mux44~16_combout ;
wire \reg_file_nxt[31][17]~87_combout ;
wire \reg_file[29][17]~q ;
wire \reg_file[17][17]~q ;
wire \reg_file[25][17]~feeder_combout ;
wire \reg_file[25][17]~q ;
wire \Mux46~0_combout ;
wire \reg_file[21][17]~feeder_combout ;
wire \reg_file[21][17]~q ;
wire \Mux46~1_combout ;
wire \reg_file[23][17]~feeder_combout ;
wire \reg_file[23][17]~q ;
wire \reg_file[31][17]~q ;
wire \reg_file[27][17]~q ;
wire \reg_file[19][17]~q ;
wire \Mux46~7_combout ;
wire \Mux46~8_combout ;
wire \reg_file[30][17]~q ;
wire \reg_file[22][17]~q ;
wire \reg_file[18][17]~q ;
wire \Mux46~2_combout ;
wire \Mux46~3_combout ;
wire \reg_file[24][17]~q ;
wire \reg_file[28][17]~q ;
wire \Mux46~5_combout ;
wire \Mux46~6_combout ;
wire \reg_file[9][17]~feeder_combout ;
wire \reg_file[9][17]~q ;
wire \reg_file[10][17]~q ;
wire \reg_file[8][17]~q ;
wire \Mux46~12_combout ;
wire \Mux46~13_combout ;
wire \reg_file[1][17]~q ;
wire \reg_file[3][17]~feeder_combout ;
wire \reg_file[3][17]~q ;
wire \Mux46~14_combout ;
wire \Mux46~15_combout ;
wire \Mux46~16_combout ;
wire \reg_file[13][17]~q ;
wire \reg_file[12][17]~q ;
wire \Mux46~17_combout ;
wire \reg_file[14][17]~q ;
wire \reg_file[15][17]~q ;
wire \Mux46~18_combout ;
wire \reg_file[7][17]~q ;
wire \reg_file[6][17]~q ;
wire \reg_file[5][17]~q ;
wire \reg_file[4][17]~q ;
wire \Mux46~10_combout ;
wire \Mux46~11_combout ;
wire \reg_file_nxt[31][21]~88_combout ;
wire \reg_file[31][21]~feeder_combout ;
wire \reg_file[31][21]~q ;
wire \reg_file[23][21]~q ;
wire \reg_file[27][21]~q ;
wire \Mux42~7_combout ;
wire \Mux42~8_combout ;
wire \reg_file[21][21]~q ;
wire \reg_file[29][21]~q ;
wire \reg_file[17][21]~q ;
wire \reg_file[25][21]~feeder_combout ;
wire \reg_file[25][21]~q ;
wire \Mux42~0_combout ;
wire \Mux42~1_combout ;
wire \reg_file[30][21]~feeder_combout ;
wire \reg_file[30][21]~q ;
wire \reg_file[26][21]~q ;
wire \reg_file[22][21]~q ;
wire \reg_file[18][21]~q ;
wire \Mux42~2_combout ;
wire \Mux42~3_combout ;
wire \reg_file[28][21]~q ;
wire \reg_file[20][21]~feeder_combout ;
wire \reg_file[20][21]~q ;
wire \reg_file[16][21]~q ;
wire \Mux42~4_combout ;
wire \Mux42~5_combout ;
wire \Mux42~6_combout ;
wire \reg_file[15][21]~q ;
wire \reg_file[14][21]~q ;
wire \reg_file[13][21]~q ;
wire \reg_file[12][21]~q ;
wire \Mux42~17_combout ;
wire \Mux42~18_combout ;
wire \reg_file[4][21]~q ;
wire \reg_file[5][21]~q ;
wire \Mux42~10_combout ;
wire \reg_file[6][21]~feeder_combout ;
wire \reg_file[6][21]~q ;
wire \reg_file[7][21]~q ;
wire \Mux42~11_combout ;
wire \reg_file[1][21]~q ;
wire \reg_file[3][21]~feeder_combout ;
wire \reg_file[3][21]~q ;
wire \Mux42~14_combout ;
wire \reg_file[2][21]~q ;
wire \Mux42~15_combout ;
wire \reg_file[11][21]~q ;
wire \reg_file[8][21]~q ;
wire \reg_file[10][21]~q ;
wire \Mux42~12_combout ;
wire \Mux42~13_combout ;
wire \Mux42~16_combout ;
wire \reg_file_nxt[31][20]~89_combout ;
wire \reg_file[27][20]~feeder_combout ;
wire \reg_file[27][20]~q ;
wire \reg_file[31][20]~q ;
wire \reg_file[23][20]~q ;
wire \reg_file[19][20]~q ;
wire \Mux43~7_combout ;
wire \Mux43~8_combout ;
wire \reg_file[29][20]~feeder_combout ;
wire \reg_file[29][20]~q ;
wire \reg_file[21][20]~q ;
wire \reg_file[17][20]~q ;
wire \Mux43~0_combout ;
wire \reg_file[25][20]~q ;
wire \Mux43~1_combout ;
wire \reg_file[20][20]~q ;
wire \reg_file[28][20]~q ;
wire \reg_file[24][20]~feeder_combout ;
wire \reg_file[24][20]~q ;
wire \reg_file[16][20]~q ;
wire \Mux43~4_combout ;
wire \Mux43~5_combout ;
wire \reg_file[22][20]~q ;
wire \reg_file[30][20]~q ;
wire \Mux43~3_combout ;
wire \Mux43~6_combout ;
wire \reg_file[11][20]~q ;
wire \reg_file[9][20]~feeder_combout ;
wire \reg_file[9][20]~q ;
wire \reg_file[10][20]~q ;
wire \Mux43~10_combout ;
wire \Mux43~11_combout ;
wire \reg_file[15][20]~q ;
wire \reg_file[14][20]~q ;
wire \reg_file[13][20]~q ;
wire \Mux43~17_combout ;
wire \Mux43~18_combout ;
wire \reg_file[5][20]~q ;
wire \reg_file[4][20]~q ;
wire \Mux43~12_combout ;
wire \reg_file[7][20]~q ;
wire \Mux43~13_combout ;
wire \reg_file[2][20]~q ;
wire \reg_file[3][20]~q ;
wire \reg_file[1][20]~feeder_combout ;
wire \reg_file[1][20]~q ;
wire \Mux43~14_combout ;
wire \Mux43~15_combout ;
wire \Mux43~16_combout ;
wire \reg_file_nxt[31][28]~90_combout ;
wire \reg_file[29][28]~feeder_combout ;
wire \reg_file[29][28]~q ;
wire \reg_file[17][28]~feeder_combout ;
wire \reg_file[17][28]~q ;
wire \reg_file[21][28]~q ;
wire \Mux35~0_combout ;
wire \reg_file[25][28]~feeder_combout ;
wire \reg_file[25][28]~q ;
wire \Mux35~1_combout ;
wire \reg_file[30][28]~q ;
wire \reg_file[22][28]~feeder_combout ;
wire \reg_file[22][28]~q ;
wire \Mux35~3_combout ;
wire \reg_file[28][28]~q ;
wire \reg_file[20][28]~q ;
wire \reg_file[24][28]~feeder_combout ;
wire \reg_file[24][28]~q ;
wire \reg_file[16][28]~q ;
wire \Mux35~4_combout ;
wire \Mux35~5_combout ;
wire \Mux35~6_combout ;
wire \reg_file[23][28]~q ;
wire \reg_file[19][28]~q ;
wire \Mux35~7_combout ;
wire \reg_file[27][28]~q ;
wire \reg_file[31][28]~q ;
wire \Mux35~8_combout ;
wire \reg_file[9][28]~feeder_combout ;
wire \reg_file[9][28]~q ;
wire \reg_file[11][28]~feeder_combout ;
wire \reg_file[11][28]~q ;
wire \reg_file[10][28]~q ;
wire \Mux35~10_combout ;
wire \Mux35~11_combout ;
wire \reg_file[14][28]~feeder_combout ;
wire \reg_file[14][28]~q ;
wire \reg_file[13][28]~q ;
wire \Mux35~17_combout ;
wire \reg_file[15][28]~q ;
wire \Mux35~18_combout ;
wire \reg_file[2][28]~feeder_combout ;
wire \reg_file[2][28]~q ;
wire \reg_file[1][28]~feeder_combout ;
wire \reg_file[1][28]~q ;
wire \reg_file[3][28]~q ;
wire \Mux35~14_combout ;
wire \Mux35~15_combout ;
wire \reg_file[7][28]~feeder_combout ;
wire \reg_file[7][28]~q ;
wire \reg_file[6][28]~q ;
wire \Mux35~13_combout ;
wire \Mux35~16_combout ;
wire \reg_file_nxt[31][26]~91_combout ;
wire \reg_file[22][26]~feeder_combout ;
wire \reg_file[22][26]~q ;
wire \reg_file[30][26]~q ;
wire \Mux37~3_combout ;
wire \reg_file[20][26]~q ;
wire \reg_file[28][26]~q ;
wire \Mux37~5_combout ;
wire \Mux37~6_combout ;
wire \reg_file[29][26]~feeder_combout ;
wire \reg_file[29][26]~q ;
wire \reg_file[25][26]~q ;
wire \reg_file[17][26]~q ;
wire \reg_file[21][26]~q ;
wire \Mux37~0_combout ;
wire \Mux37~1_combout ;
wire \reg_file[31][26]~q ;
wire \reg_file[27][26]~q ;
wire \reg_file[23][26]~q ;
wire \reg_file[19][26]~q ;
wire \Mux37~7_combout ;
wire \Mux37~8_combout ;
wire \reg_file[10][26]~q ;
wire \Mux37~10_combout ;
wire \reg_file[9][26]~q ;
wire \reg_file[11][26]~feeder_combout ;
wire \reg_file[11][26]~q ;
wire \Mux37~11_combout ;
wire \reg_file[15][26]~q ;
wire \reg_file[14][26]~q ;
wire \reg_file[13][26]~q ;
wire \Mux37~17_combout ;
wire \Mux37~18_combout ;
wire \reg_file[6][26]~q ;
wire \reg_file[7][26]~q ;
wire \reg_file[5][26]~q ;
wire \Mux37~12_combout ;
wire \Mux37~13_combout ;
wire \reg_file[1][26]~q ;
wire \reg_file[3][26]~q ;
wire \Mux37~14_combout ;
wire \reg_file[2][26]~q ;
wire \Mux37~15_combout ;
wire \Mux37~16_combout ;
wire \reg_file_nxt[31][8]~92_combout ;
wire \reg_file[29][8]~q ;
wire \reg_file[17][8]~q ;
wire \Mux55~0_combout ;
wire \reg_file[25][8]~feeder_combout ;
wire \reg_file[25][8]~q ;
wire \Mux55~1_combout ;
wire \reg_file[23][8]~q ;
wire \reg_file[19][8]~q ;
wire \Mux55~7_combout ;
wire \reg_file[27][8]~q ;
wire \reg_file[31][8]~feeder_combout ;
wire \reg_file[31][8]~q ;
wire \Mux55~8_combout ;
wire \reg_file[20][8]~q ;
wire \reg_file[28][8]~q ;
wire \reg_file[16][8]~q ;
wire \reg_file[24][8]~feeder_combout ;
wire \reg_file[24][8]~q ;
wire \Mux55~4_combout ;
wire \Mux55~5_combout ;
wire \reg_file[18][8]~q ;
wire \reg_file[26][8]~q ;
wire \Mux55~2_combout ;
wire \reg_file[22][8]~q ;
wire \Mux55~3_combout ;
wire \Mux55~6_combout ;
wire \reg_file[2][8]~feeder_combout ;
wire \reg_file[2][8]~q ;
wire \reg_file[1][8]~q ;
wire \reg_file[3][8]~q ;
wire \Mux55~14_combout ;
wire \Mux55~15_combout ;
wire \reg_file[6][8]~q ;
wire \reg_file[5][8]~q ;
wire \reg_file[4][8]~q ;
wire \Mux55~12_combout ;
wire \Mux55~13_combout ;
wire \Mux55~16_combout ;
wire \reg_file[8][8]~q ;
wire \reg_file[10][8]~q ;
wire \Mux55~10_combout ;
wire \reg_file[11][8]~q ;
wire \reg_file[9][8]~q ;
wire \Mux55~11_combout ;
wire \reg_file[15][8]~feeder_combout ;
wire \reg_file[15][8]~q ;
wire \reg_file[14][8]~q ;
wire \reg_file[12][8]~q ;
wire \reg_file[13][8]~q ;
wire \Mux55~17_combout ;
wire \Mux55~18_combout ;
wire \reg_file_nxt[31][7]~93_combout ;
wire \reg_file[19][7]~q ;
wire \reg_file[27][7]~q ;
wire \Mux56~7_combout ;
wire \reg_file[23][7]~feeder_combout ;
wire \reg_file[23][7]~q ;
wire \reg_file[31][7]~q ;
wire \Mux56~8_combout ;
wire \reg_file[29][7]~feeder_combout ;
wire \reg_file[29][7]~q ;
wire \reg_file[21][7]~feeder_combout ;
wire \reg_file[21][7]~q ;
wire \reg_file[17][7]~feeder_combout ;
wire \reg_file[17][7]~q ;
wire \reg_file[25][7]~q ;
wire \Mux56~0_combout ;
wire \Mux56~1_combout ;
wire \reg_file[24][7]~q ;
wire \reg_file[20][7]~feeder_combout ;
wire \reg_file[20][7]~q ;
wire \Mux56~4_combout ;
wire \reg_file[28][7]~q ;
wire \Mux56~5_combout ;
wire \reg_file[22][7]~q ;
wire \Mux56~2_combout ;
wire \reg_file[26][7]~q ;
wire \reg_file[30][7]~feeder_combout ;
wire \reg_file[30][7]~q ;
wire \Mux56~3_combout ;
wire \Mux56~6_combout ;
wire \reg_file[4][7]~q ;
wire \reg_file[5][7]~q ;
wire \Mux56~10_combout ;
wire \reg_file[6][7]~q ;
wire \reg_file[7][7]~q ;
wire \Mux56~11_combout ;
wire \reg_file[12][7]~q ;
wire \reg_file[13][7]~q ;
wire \Mux56~17_combout ;
wire \reg_file[15][7]~feeder_combout ;
wire \reg_file[15][7]~q ;
wire \reg_file[14][7]~feeder_combout ;
wire \reg_file[14][7]~q ;
wire \Mux56~18_combout ;
wire \reg_file[2][7]~feeder_combout ;
wire \reg_file[2][7]~q ;
wire \reg_file[1][7]~q ;
wire \reg_file[3][7]~q ;
wire \Mux56~14_combout ;
wire \Mux56~15_combout ;
wire \reg_file[11][7]~feeder_combout ;
wire \reg_file[11][7]~q ;
wire \reg_file[8][7]~q ;
wire \reg_file[10][7]~q ;
wire \Mux56~12_combout ;
wire \Mux56~13_combout ;
wire \Mux56~16_combout ;
wire \reg_file_nxt[31][22]~94_combout ;
wire \reg_file[29][22]~feeder_combout ;
wire \reg_file[29][22]~q ;
wire \reg_file[25][22]~q ;
wire \reg_file[17][22]~q ;
wire \reg_file[21][22]~q ;
wire \Mux41~0_combout ;
wire \Mux41~1_combout ;
wire \reg_file[27][22]~feeder_combout ;
wire \reg_file[27][22]~q ;
wire \reg_file[31][22]~q ;
wire \reg_file[23][22]~q ;
wire \reg_file[19][22]~q ;
wire \Mux41~7_combout ;
wire \Mux41~8_combout ;
wire \reg_file[28][22]~q ;
wire \reg_file[20][22]~q ;
wire \reg_file[24][22]~q ;
wire \Mux41~4_combout ;
wire \Mux41~5_combout ;
wire \reg_file[22][22]~feeder_combout ;
wire \reg_file[22][22]~q ;
wire \reg_file[30][22]~q ;
wire \reg_file[18][22]~q ;
wire \reg_file[26][22]~q ;
wire \Mux41~2_combout ;
wire \Mux41~3_combout ;
wire \Mux41~6_combout ;
wire \reg_file[13][22]~q ;
wire \reg_file[12][22]~q ;
wire \Mux41~17_combout ;
wire \reg_file[14][22]~q ;
wire \reg_file[15][22]~q ;
wire \Mux41~18_combout ;
wire \reg_file[11][22]~q ;
wire \reg_file[9][22]~q ;
wire \reg_file[8][22]~q ;
wire \reg_file[10][22]~q ;
wire \Mux41~10_combout ;
wire \Mux41~11_combout ;
wire \reg_file[3][22]~q ;
wire \reg_file[1][22]~q ;
wire \Mux41~14_combout ;
wire \reg_file[2][22]~q ;
wire \Mux41~15_combout ;
wire \reg_file[7][22]~feeder_combout ;
wire \reg_file[7][22]~q ;
wire \reg_file[5][22]~q ;
wire \reg_file[4][22]~q ;
wire \Mux41~12_combout ;
wire \reg_file[6][22]~q ;
wire \Mux41~13_combout ;
wire \Mux41~16_combout ;
wire \reg_file_nxt[31][25]~95_combout ;
wire \reg_file[23][25]~feeder_combout ;
wire \reg_file[23][25]~q ;
wire \reg_file[27][25]~q ;
wire \reg_file[19][25]~q ;
wire \Mux38~7_combout ;
wire \reg_file[31][25]~q ;
wire \Mux38~8_combout ;
wire \reg_file[25][25]~q ;
wire \reg_file[17][25]~feeder_combout ;
wire \reg_file[17][25]~q ;
wire \Mux38~0_combout ;
wire \reg_file[21][25]~q ;
wire \reg_file[29][25]~feeder_combout ;
wire \reg_file[29][25]~q ;
wire \Mux38~1_combout ;
wire \reg_file[28][25]~q ;
wire \reg_file[24][25]~q ;
wire \Mux38~5_combout ;
wire \reg_file[18][25]~feeder_combout ;
wire \reg_file[18][25]~q ;
wire \reg_file[22][25]~feeder_combout ;
wire \reg_file[22][25]~q ;
wire \Mux38~2_combout ;
wire \reg_file[30][25]~q ;
wire \reg_file[26][25]~feeder_combout ;
wire \reg_file[26][25]~q ;
wire \Mux38~3_combout ;
wire \Mux38~6_combout ;
wire \reg_file[15][25]~q ;
wire \reg_file[14][25]~q ;
wire \reg_file[13][25]~q ;
wire \reg_file[12][25]~q ;
wire \Mux38~17_combout ;
wire \Mux38~18_combout ;
wire \reg_file[2][25]~q ;
wire \Mux38~15_combout ;
wire \reg_file[9][25]~q ;
wire \reg_file[11][25]~q ;
wire \reg_file[8][25]~q ;
wire \reg_file[10][25]~q ;
wire \Mux38~12_combout ;
wire \Mux38~13_combout ;
wire \Mux38~16_combout ;
wire \reg_file[7][25]~q ;
wire \reg_file[6][25]~q ;
wire \reg_file[5][25]~q ;
wire \reg_file[4][25]~q ;
wire \Mux38~10_combout ;
wire \Mux38~11_combout ;
wire \Mux29~0_combout ;
wire \Mux29~1_combout ;
wire \Mux29~7_combout ;
wire \Mux29~8_combout ;
wire \reg_file[28][2]~q ;
wire \Mux29~5_combout ;
wire \Mux29~2_combout ;
wire \reg_file[30][2]~q ;
wire \Mux29~3_combout ;
wire \Mux29~6_combout ;
wire \Mux29~17_combout ;
wire \Mux29~18_combout ;
wire \reg_file[6][2]~q ;
wire \Mux29~10_combout ;
wire \Mux29~11_combout ;
wire \Mux29~15_combout ;
wire \Mux29~13_combout ;
wire \Mux29~16_combout ;
wire \Mux27~0_combout ;
wire \Mux27~1_combout ;
wire \Mux27~7_combout ;
wire \Mux27~8_combout ;
wire \reg_file[16][4]~q ;
wire \Mux27~4_combout ;
wire \reg_file[24][4]~q ;
wire \Mux27~5_combout ;
wire \Mux27~3_combout ;
wire \Mux27~6_combout ;
wire \reg_file[6][4]~feeder_combout ;
wire \reg_file[6][4]~q ;
wire \Mux27~10_combout ;
wire \Mux27~11_combout ;
wire \Mux27~17_combout ;
wire \Mux27~18_combout ;
wire \reg_file[3][4]~q ;
wire \Mux27~14_combout ;
wire \Mux27~15_combout ;
wire \Mux27~13_combout ;
wire \Mux27~16_combout ;
wire \Mux28~7_combout ;
wire \Mux28~8_combout ;
wire \reg_file[26][3]~q ;
wire \Mux28~2_combout ;
wire \Mux28~3_combout ;
wire \reg_file[24][3]~q ;
wire \Mux28~4_combout ;
wire \Mux28~5_combout ;
wire \Mux28~6_combout ;
wire \Mux28~0_combout ;
wire \Mux28~1_combout ;
wire \Mux28~15_combout ;
wire \Mux28~12_combout ;
wire \Mux28~13_combout ;
wire \Mux28~16_combout ;
wire \Mux28~10_combout ;
wire \Mux28~11_combout ;
wire \Mux28~17_combout ;
wire \Mux28~18_combout ;
wire \Mux23~7_combout ;
wire \Mux23~8_combout ;
wire \Mux23~2_combout ;
wire \reg_file[30][8]~q ;
wire \Mux23~3_combout ;
wire \Mux23~4_combout ;
wire \Mux23~5_combout ;
wire \Mux23~6_combout ;
wire \reg_file[21][8]~feeder_combout ;
wire \reg_file[21][8]~q ;
wire \Mux23~0_combout ;
wire \Mux23~1_combout ;
wire \Mux23~10_combout ;
wire \reg_file[7][8]~feeder_combout ;
wire \reg_file[7][8]~q ;
wire \Mux23~11_combout ;
wire \Mux23~17_combout ;
wire \Mux23~18_combout ;
wire \Mux23~15_combout ;
wire \Mux23~12_combout ;
wire \Mux23~13_combout ;
wire \Mux23~16_combout ;
wire \Mux24~7_combout ;
wire \Mux24~8_combout ;
wire \reg_file[16][7]~feeder_combout ;
wire \reg_file[16][7]~q ;
wire \Mux24~4_combout ;
wire \Mux24~5_combout ;
wire \reg_file[18][7]~q ;
wire \Mux24~2_combout ;
wire \Mux24~3_combout ;
wire \Mux24~6_combout ;
wire \Mux24~0_combout ;
wire \Mux24~1_combout ;
wire \Mux24~17_combout ;
wire \Mux24~18_combout ;
wire \Mux24~10_combout ;
wire \reg_file[9][7]~q ;
wire \Mux24~11_combout ;
wire \Mux24~12_combout ;
wire \Mux24~13_combout ;
wire \Mux24~14_combout ;
wire \Mux24~15_combout ;
wire \Mux24~16_combout ;
wire \Mux25~7_combout ;
wire \Mux25~8_combout ;
wire \reg_file[20][6]~q ;
wire \Mux25~4_combout ;
wire \Mux25~5_combout ;
wire \reg_file[30][6]~q ;
wire \Mux25~3_combout ;
wire \Mux25~6_combout ;
wire \reg_file[21][6]~q ;
wire \Mux25~0_combout ;
wire \Mux25~1_combout ;
wire \Mux25~17_combout ;
wire \Mux25~18_combout ;
wire \Mux25~12_combout ;
wire \Mux25~13_combout ;
wire \Mux25~14_combout ;
wire \Mux25~15_combout ;
wire \Mux25~16_combout ;
wire \Mux25~10_combout ;
wire \Mux25~11_combout ;
wire \Mux26~0_combout ;
wire \Mux26~1_combout ;
wire \Mux26~7_combout ;
wire \Mux26~8_combout ;
wire \Mux26~4_combout ;
wire \reg_file[28][5]~q ;
wire \Mux26~5_combout ;
wire \reg_file[22][5]~feeder_combout ;
wire \reg_file[22][5]~q ;
wire \reg_file[18][5]~q ;
wire \Mux26~2_combout ;
wire \Mux26~3_combout ;
wire \Mux26~6_combout ;
wire \reg_file[2][5]~feeder_combout ;
wire \reg_file[2][5]~q ;
wire \Mux26~14_combout ;
wire \Mux26~15_combout ;
wire \Mux26~12_combout ;
wire \Mux26~13_combout ;
wire \Mux26~16_combout ;
wire \Mux26~17_combout ;
wire \Mux26~18_combout ;
wire \Mux26~10_combout ;
wire \Mux26~11_combout ;
wire \reg_file[19][16]~q ;
wire \Mux15~7_combout ;
wire \Mux15~8_combout ;
wire \reg_file[21][16]~feeder_combout ;
wire \reg_file[21][16]~q ;
wire \Mux15~0_combout ;
wire \Mux15~1_combout ;
wire \reg_file[26][16]~q ;
wire \reg_file[18][16]~q ;
wire \Mux15~2_combout ;
wire \Mux15~3_combout ;
wire \Mux15~4_combout ;
wire \Mux15~5_combout ;
wire \Mux15~6_combout ;
wire \Mux15~17_combout ;
wire \Mux15~18_combout ;
wire \Mux15~13_combout ;
wire \reg_file[3][16]~feeder_combout ;
wire \reg_file[3][16]~q ;
wire \Mux15~14_combout ;
wire \Mux15~15_combout ;
wire \Mux15~16_combout ;
wire \Mux15~10_combout ;
wire \Mux15~11_combout ;
wire \Mux16~0_combout ;
wire \Mux16~1_combout ;
wire \Mux16~7_combout ;
wire \Mux16~8_combout ;
wire \Mux16~2_combout ;
wire \Mux16~3_combout ;
wire \Mux16~4_combout ;
wire \Mux16~5_combout ;
wire \Mux16~6_combout ;
wire \Mux16~17_combout ;
wire \Mux16~18_combout ;
wire \Mux16~10_combout ;
wire \Mux16~11_combout ;
wire \Mux16~14_combout ;
wire \Mux16~15_combout ;
wire \Mux16~12_combout ;
wire \Mux16~13_combout ;
wire \Mux16~16_combout ;
wire \Mux17~0_combout ;
wire \Mux17~1_combout ;
wire \Mux17~7_combout ;
wire \Mux17~8_combout ;
wire \Mux17~4_combout ;
wire \Mux17~5_combout ;
wire \reg_file[30][14]~feeder_combout ;
wire \reg_file[30][14]~q ;
wire \Mux17~2_combout ;
wire \Mux17~3_combout ;
wire \Mux17~6_combout ;
wire \Mux17~15_combout ;
wire \reg_file[8][14]~q ;
wire \Mux17~12_combout ;
wire \Mux17~13_combout ;
wire \Mux17~16_combout ;
wire \Mux17~17_combout ;
wire \Mux17~18_combout ;
wire \Mux17~10_combout ;
wire \Mux17~11_combout ;
wire \reg_file[17][13]~feeder_combout ;
wire \reg_file[17][13]~q ;
wire \Mux18~0_combout ;
wire \Mux18~1_combout ;
wire \Mux18~7_combout ;
wire \Mux18~8_combout ;
wire \reg_file[26][13]~q ;
wire \Mux18~2_combout ;
wire \Mux18~3_combout ;
wire \reg_file[28][13]~q ;
wire \reg_file[16][13]~q ;
wire \Mux18~4_combout ;
wire \Mux18~5_combout ;
wire \Mux18~6_combout ;
wire \reg_file[12][13]~q ;
wire \Mux18~17_combout ;
wire \Mux18~18_combout ;
wire \reg_file[8][13]~q ;
wire \reg_file[10][13]~q ;
wire \Mux18~10_combout ;
wire \Mux18~11_combout ;
wire \Mux18~14_combout ;
wire \Mux18~15_combout ;
wire \Mux18~13_combout ;
wire \Mux18~16_combout ;
wire \Mux20~2_combout ;
wire \Mux20~3_combout ;
wire \Mux20~4_combout ;
wire \Mux20~5_combout ;
wire \Mux20~6_combout ;
wire \reg_file[17][11]~q ;
wire \Mux20~0_combout ;
wire \Mux20~1_combout ;
wire \Mux20~7_combout ;
wire \Mux20~8_combout ;
wire \Mux20~12_combout ;
wire \Mux20~13_combout ;
wire \Mux20~14_combout ;
wire \Mux20~15_combout ;
wire \Mux20~16_combout ;
wire \reg_file[8][11]~q ;
wire \reg_file[10][11]~q ;
wire \Mux20~10_combout ;
wire \Mux20~11_combout ;
wire \Mux20~17_combout ;
wire \Mux20~18_combout ;
wire \Mux19~7_combout ;
wire \Mux19~8_combout ;
wire \Mux19~0_combout ;
wire \Mux19~1_combout ;
wire \Mux19~3_combout ;
wire \Mux19~4_combout ;
wire \Mux19~5_combout ;
wire \Mux19~6_combout ;
wire \reg_file[6][12]~feeder_combout ;
wire \reg_file[6][12]~q ;
wire \Mux19~10_combout ;
wire \Mux19~11_combout ;
wire \Mux19~17_combout ;
wire \Mux19~18_combout ;
wire \Mux19~13_combout ;
wire \Mux19~15_combout ;
wire \Mux19~16_combout ;
wire \Mux21~7_combout ;
wire \Mux21~8_combout ;
wire \Mux21~2_combout ;
wire \Mux21~3_combout ;
wire \Mux21~4_combout ;
wire \reg_file[28][10]~q ;
wire \Mux21~5_combout ;
wire \Mux21~6_combout ;
wire \Mux21~0_combout ;
wire \Mux21~1_combout ;
wire \Mux21~10_combout ;
wire \Mux21~11_combout ;
wire \Mux21~17_combout ;
wire \Mux21~18_combout ;
wire \Mux21~14_combout ;
wire \Mux21~15_combout ;
wire \Mux21~13_combout ;
wire \Mux21~16_combout ;
wire \Mux22~0_combout ;
wire \Mux22~1_combout ;
wire \reg_file[19][9]~q ;
wire \Mux22~7_combout ;
wire \Mux22~8_combout ;
wire \Mux22~4_combout ;
wire \Mux22~5_combout ;
wire \Mux22~3_combout ;
wire \Mux22~6_combout ;
wire \Mux22~17_combout ;
wire \Mux22~18_combout ;
wire \reg_file[10][9]~q ;
wire \reg_file[8][9]~q ;
wire \Mux22~10_combout ;
wire \Mux22~11_combout ;
wire \Mux22~15_combout ;
wire \Mux22~12_combout ;
wire \Mux22~13_combout ;
wire \Mux22~16_combout ;
wire \Mux13~7_combout ;
wire \Mux13~8_combout ;
wire \Mux13~0_combout ;
wire \Mux13~1_combout ;
wire \Mux13~2_combout ;
wire \Mux13~3_combout ;
wire \reg_file[24][18]~feeder_combout ;
wire \reg_file[24][18]~q ;
wire \Mux13~5_combout ;
wire \Mux13~6_combout ;
wire \reg_file[4][18]~q ;
wire \reg_file[5][18]~q ;
wire \Mux13~10_combout ;
wire \Mux13~11_combout ;
wire \reg_file[12][18]~q ;
wire \Mux13~17_combout ;
wire \Mux13~18_combout ;
wire \reg_file[3][18]~q ;
wire \Mux13~14_combout ;
wire \Mux13~15_combout ;
wire \Mux13~13_combout ;
wire \Mux13~16_combout ;
wire \Mux14~0_combout ;
wire \Mux14~1_combout ;
wire \reg_file[26][17]~feeder_combout ;
wire \reg_file[26][17]~q ;
wire \Mux14~2_combout ;
wire \Mux14~3_combout ;
wire \reg_file[16][17]~q ;
wire \Mux14~4_combout ;
wire \Mux14~5_combout ;
wire \Mux14~6_combout ;
wire \Mux14~7_combout ;
wire \Mux14~8_combout ;
wire \Mux14~17_combout ;
wire \Mux14~18_combout ;
wire \reg_file[2][17]~q ;
wire \Mux14~15_combout ;
wire \Mux14~13_combout ;
wire \Mux14~16_combout ;
wire \Mux14~10_combout ;
wire \reg_file[11][17]~q ;
wire \Mux14~11_combout ;
wire \Mux11~0_combout ;
wire \Mux11~1_combout ;
wire \Mux11~7_combout ;
wire \Mux11~8_combout ;
wire \reg_file[26][20]~q ;
wire \reg_file[18][20]~q ;
wire \Mux11~2_combout ;
wire \Mux11~3_combout ;
wire \Mux11~4_combout ;
wire \Mux11~5_combout ;
wire \Mux11~6_combout ;
wire \reg_file[12][20]~q ;
wire \Mux11~17_combout ;
wire \Mux11~18_combout ;
wire \reg_file[6][20]~feeder_combout ;
wire \reg_file[6][20]~q ;
wire \Mux11~10_combout ;
wire \Mux11~11_combout ;
wire \Mux11~13_combout ;
wire \Mux11~15_combout ;
wire \Mux11~16_combout ;
wire \Mux12~0_combout ;
wire \Mux12~1_combout ;
wire \Mux12~3_combout ;
wire \reg_file[24][19]~q ;
wire \Mux12~4_combout ;
wire \Mux12~5_combout ;
wire \Mux12~6_combout ;
wire \Mux12~7_combout ;
wire \Mux12~8_combout ;
wire \reg_file[11][19]~feeder_combout ;
wire \reg_file[11][19]~q ;
wire \Mux12~10_combout ;
wire \Mux12~11_combout ;
wire \Mux12~17_combout ;
wire \Mux12~18_combout ;
wire \Mux12~12_combout ;
wire \Mux12~13_combout ;
wire \Mux12~14_combout ;
wire \Mux12~15_combout ;
wire \Mux12~16_combout ;
wire \Mux9~0_combout ;
wire \Mux9~1_combout ;
wire \Mux9~7_combout ;
wire \Mux9~8_combout ;
wire \Mux9~2_combout ;
wire \Mux9~3_combout ;
wire \reg_file[16][22]~q ;
wire \Mux9~4_combout ;
wire \Mux9~5_combout ;
wire \Mux9~6_combout ;
wire \Mux9~17_combout ;
wire \Mux9~18_combout ;
wire \Mux9~10_combout ;
wire \Mux9~11_combout ;
wire \Mux9~12_combout ;
wire \Mux9~13_combout ;
wire \Mux9~14_combout ;
wire \Mux9~15_combout ;
wire \Mux9~16_combout ;
wire \reg_file[24][21]~q ;
wire \Mux10~4_combout ;
wire \Mux10~5_combout ;
wire \Mux10~2_combout ;
wire \Mux10~3_combout ;
wire \Mux10~6_combout ;
wire \reg_file[19][21]~q ;
wire \Mux10~7_combout ;
wire \Mux10~8_combout ;
wire \Mux10~0_combout ;
wire \Mux10~1_combout ;
wire \Mux10~10_combout ;
wire \reg_file[9][21]~q ;
wire \Mux10~11_combout ;
wire \Mux10~17_combout ;
wire \Mux10~18_combout ;
wire \Mux10~12_combout ;
wire \Mux10~13_combout ;
wire \Mux10~14_combout ;
wire \Mux10~15_combout ;
wire \Mux10~16_combout ;
wire \Mux7~7_combout ;
wire \Mux7~8_combout ;
wire \Mux7~0_combout ;
wire \Mux7~1_combout ;
wire \reg_file[30][24]~feeder_combout ;
wire \reg_file[30][24]~q ;
wire \Mux7~3_combout ;
wire \reg_file[24][24]~feeder_combout ;
wire \reg_file[24][24]~q ;
wire \Mux7~5_combout ;
wire \Mux7~6_combout ;
wire \Mux7~17_combout ;
wire \Mux7~18_combout ;
wire \Mux7~10_combout ;
wire \Mux7~11_combout ;
wire \Mux7~13_combout ;
wire \Mux7~15_combout ;
wire \Mux7~16_combout ;
wire \Mux8~2_combout ;
wire \Mux8~3_combout ;
wire \reg_file[20][23]~q ;
wire \reg_file[16][23]~q ;
wire \Mux8~4_combout ;
wire \Mux8~5_combout ;
wire \Mux8~6_combout ;
wire \reg_file[17][23]~feeder_combout ;
wire \reg_file[17][23]~q ;
wire \Mux8~0_combout ;
wire \Mux8~1_combout ;
wire \Mux8~7_combout ;
wire \Mux8~8_combout ;
wire \Mux8~14_combout ;
wire \Mux8~15_combout ;
wire \Mux8~12_combout ;
wire \Mux8~13_combout ;
wire \Mux8~16_combout ;
wire \reg_file[9][23]~q ;
wire \Mux8~10_combout ;
wire \Mux8~11_combout ;
wire \Mux8~17_combout ;
wire \Mux8~18_combout ;
wire \Mux0~0_combout ;
wire \Mux0~1_combout ;
wire \Mux0~7_combout ;
wire \Mux0~8_combout ;
wire \reg_file[22][31]~q ;
wire \Mux0~3_combout ;
wire \reg_file[20][31]~q ;
wire \reg_file[16][31]~q ;
wire \Mux0~4_combout ;
wire \Mux0~5_combout ;
wire \Mux0~6_combout ;
wire \Mux0~17_combout ;
wire \Mux0~18_combout ;
wire \Mux0~10_combout ;
wire \Mux0~11_combout ;
wire \Mux0~12_combout ;
wire \Mux0~13_combout ;
wire \Mux0~14_combout ;
wire \Mux0~15_combout ;
wire \Mux0~16_combout ;
wire \Mux1~0_combout ;
wire \Mux1~1_combout ;
wire \Mux1~7_combout ;
wire \Mux1~8_combout ;
wire \Mux1~3_combout ;
wire \reg_file[24][30]~q ;
wire \reg_file[16][30]~q ;
wire \Mux1~4_combout ;
wire \Mux1~5_combout ;
wire \Mux1~6_combout ;
wire \Mux1~17_combout ;
wire \Mux1~18_combout ;
wire \reg_file[7][30]~feeder_combout ;
wire \reg_file[7][30]~q ;
wire \Mux1~10_combout ;
wire \Mux1~11_combout ;
wire \Mux1~13_combout ;
wire \reg_file[1][30]~q ;
wire \reg_file[3][30]~q ;
wire \Mux1~14_combout ;
wire \Mux1~15_combout ;
wire \Mux1~16_combout ;
wire \Mux2~3_combout ;
wire \reg_file[20][29]~feeder_combout ;
wire \reg_file[20][29]~q ;
wire \reg_file[16][29]~q ;
wire \Mux2~4_combout ;
wire \Mux2~5_combout ;
wire \Mux2~6_combout ;
wire \Mux2~0_combout ;
wire \Mux2~1_combout ;
wire \Mux2~7_combout ;
wire \Mux2~8_combout ;
wire \Mux2~12_combout ;
wire \Mux2~13_combout ;
wire \Mux2~14_combout ;
wire \Mux2~15_combout ;
wire \Mux2~16_combout ;
wire \Mux2~17_combout ;
wire \Mux2~18_combout ;
wire \reg_file[9][29]~q ;
wire \Mux2~10_combout ;
wire \Mux2~11_combout ;
wire \Mux5~7_combout ;
wire \Mux5~8_combout ;
wire \Mux5~0_combout ;
wire \Mux5~1_combout ;
wire \reg_file[16][26]~q ;
wire \Mux5~4_combout ;
wire \Mux5~5_combout ;
wire \reg_file[18][26]~q ;
wire \Mux5~2_combout ;
wire \reg_file[26][26]~q ;
wire \Mux5~3_combout ;
wire \Mux5~6_combout ;
wire \reg_file[12][26]~q ;
wire \Mux5~17_combout ;
wire \Mux5~18_combout ;
wire \reg_file[4][26]~q ;
wire \Mux5~10_combout ;
wire \Mux5~11_combout ;
wire \Mux5~14_combout ;
wire \Mux5~15_combout ;
wire \reg_file[8][26]~q ;
wire \Mux5~12_combout ;
wire \Mux5~13_combout ;
wire \Mux5~16_combout ;
wire \Mux6~0_combout ;
wire \Mux6~1_combout ;
wire \Mux6~7_combout ;
wire \Mux6~8_combout ;
wire \reg_file[20][25]~q ;
wire \reg_file[16][25]~q ;
wire \Mux6~4_combout ;
wire \Mux6~5_combout ;
wire \Mux6~3_combout ;
wire \Mux6~6_combout ;
wire \Mux6~10_combout ;
wire \Mux6~11_combout ;
wire \reg_file[3][25]~q ;
wire \reg_file[1][25]~q ;
wire \Mux6~14_combout ;
wire \Mux6~15_combout ;
wire \Mux6~12_combout ;
wire \Mux6~13_combout ;
wire \Mux6~16_combout ;
wire \Mux6~17_combout ;
wire \Mux6~18_combout ;
wire \Mux3~7_combout ;
wire \Mux3~8_combout ;
wire \Mux3~0_combout ;
wire \Mux3~1_combout ;
wire \Mux3~5_combout ;
wire \reg_file[26][28]~q ;
wire \Mux3~3_combout ;
wire \Mux3~6_combout ;
wire \reg_file[5][28]~q ;
wire \reg_file[4][28]~q ;
wire \Mux3~10_combout ;
wire \Mux3~11_combout ;
wire \Mux3~14_combout ;
wire \Mux3~15_combout ;
wire \reg_file[8][28]~q ;
wire \Mux3~12_combout ;
wire \Mux3~13_combout ;
wire \Mux3~16_combout ;
wire \reg_file[12][28]~q ;
wire \Mux3~17_combout ;
wire \Mux3~18_combout ;
wire \Mux4~0_combout ;
wire \reg_file[25][27]~feeder_combout ;
wire \reg_file[25][27]~q ;
wire \Mux4~1_combout ;
wire \reg_file[18][27]~feeder_combout ;
wire \reg_file[18][27]~q ;
wire \Mux4~2_combout ;
wire \reg_file[22][27]~feeder_combout ;
wire \reg_file[22][27]~q ;
wire \Mux4~3_combout ;
wire \reg_file[16][27]~q ;
wire \Mux4~4_combout ;
wire \Mux4~5_combout ;
wire \Mux4~6_combout ;
wire \Mux4~7_combout ;
wire \Mux4~8_combout ;
wire \Mux4~10_combout ;
wire \Mux4~11_combout ;
wire \Mux4~14_combout ;
wire \Mux4~15_combout ;
wire \Mux4~12_combout ;
wire \Mux4~13_combout ;
wire \Mux4~16_combout ;
wire \Mux4~17_combout ;
wire \Mux4~18_combout ;


// Location: LCCOMB_X66_Y34_N2
cycloneive_lcell_comb \Mux30~4 (
// Equation(s):
// \Mux30~4_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[24][1]~q ))) # (!\prif.imemload_id [24] & (\reg_file[16][1]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][1]~q ),
	.datad(\reg_file[24][1]~q ),
	.cin(gnd),
	.combout(\Mux30~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~4 .lut_mask = 16'hDC98;
defparam \Mux30~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N4
cycloneive_lcell_comb \Mux30~14 (
// Equation(s):
// \Mux30~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][1]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][1]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[1][1]~q ),
	.datad(\reg_file[3][1]~q ),
	.cin(gnd),
	.combout(\Mux30~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~14 .lut_mask = 16'hC840;
defparam \Mux30~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y26_N23
dffeas \reg_file[4][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][0] .is_wysiwyg = "true";
defparam \reg_file[4][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N22
cycloneive_lcell_comb \Mux63~12 (
// Equation(s):
// \Mux63~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][0]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][0]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][0]~q ),
	.datad(\reg_file[5][0]~q ),
	.cin(gnd),
	.combout(\Mux63~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~12 .lut_mask = 16'hBA98;
defparam \Mux63~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N2
cycloneive_lcell_comb \Mux31~12 (
// Equation(s):
// \Mux31~12_combout  = (\prif.imemload_id [22] & ((\reg_file[10][0]~q ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\reg_file[8][0]~q  & !\prif.imemload_id [21]))))

	.dataa(\reg_file[10][0]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[8][0]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux31~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~12 .lut_mask = 16'hCCB8;
defparam \Mux31~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N31
dffeas \reg_file[16][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][2] .is_wysiwyg = "true";
defparam \reg_file[16][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N27
dffeas \reg_file[8][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][2] .is_wysiwyg = "true";
defparam \reg_file[8][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N24
cycloneive_lcell_comb \Mux59~4 (
// Equation(s):
// \Mux59~4_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[24][4]~q )) # (!\prif.imemload_id [19] & ((\reg_file[16][4]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[24][4]~q ),
	.datad(\reg_file[16][4]~q ),
	.cin(gnd),
	.combout(\Mux59~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~4 .lut_mask = 16'hD9C8;
defparam \Mux59~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y25_N31
dffeas \reg_file[8][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][4] .is_wysiwyg = "true";
defparam \reg_file[8][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N0
cycloneive_lcell_comb \Mux32~4 (
// Equation(s):
// \Mux32~4_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[20][31]~q )) # (!\prif.imemload_id [18] & ((\reg_file[16][31]~q )))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[20][31]~q ),
	.datad(\reg_file[16][31]~q ),
	.cin(gnd),
	.combout(\Mux32~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~4 .lut_mask = 16'hD9C8;
defparam \Mux32~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N26
cycloneive_lcell_comb \Mux33~4 (
// Equation(s):
// \Mux33~4_combout  = (\prif.imemload_id [19] & ((\reg_file[24][30]~q ) # ((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (((\reg_file[16][30]~q  & !\prif.imemload_id [18]))))

	.dataa(\reg_file[24][30]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[16][30]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux33~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~4 .lut_mask = 16'hCCB8;
defparam \Mux33~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N16
cycloneive_lcell_comb \Mux33~14 (
// Equation(s):
// \Mux33~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][30]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][30]~q )))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[3][30]~q ),
	.datad(\reg_file[1][30]~q ),
	.cin(gnd),
	.combout(\Mux33~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~14 .lut_mask = 16'hC480;
defparam \Mux33~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N18
cycloneive_lcell_comb \Mux34~4 (
// Equation(s):
// \Mux34~4_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[20][29]~q )) # (!\prif.imemload_id [18] & ((\reg_file[16][29]~q )))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[20][29]~q ),
	.datac(\reg_file[16][29]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux34~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~4 .lut_mask = 16'hEE50;
defparam \Mux34~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N12
cycloneive_lcell_comb \Mux58~2 (
// Equation(s):
// \Mux58~2_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[22][5]~q )) # (!\prif.imemload_id [18] & ((\reg_file[18][5]~q )))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[22][5]~q ),
	.datac(\reg_file[18][5]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux58~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~2 .lut_mask = 16'hEE50;
defparam \Mux58~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N12
cycloneive_lcell_comb \Mux50~12 (
// Equation(s):
// \Mux50~12_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][13]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][13]~q ))))

	.dataa(\reg_file[8][13]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[10][13]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux50~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~12 .lut_mask = 16'hFC22;
defparam \Mux50~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N16
cycloneive_lcell_comb \Mux52~12 (
// Equation(s):
// \Mux52~12_combout  = (\prif.imemload_id [17] & (((\reg_file[10][11]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][11]~q  & ((!\prif.imemload_id [16]))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[8][11]~q ),
	.datac(\reg_file[10][11]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux52~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~12 .lut_mask = 16'hAAE4;
defparam \Mux52~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N10
cycloneive_lcell_comb \Mux54~12 (
// Equation(s):
// \Mux54~12_combout  = (\prif.imemload_id [17] & ((\reg_file[10][9]~q ) # ((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (((\reg_file[8][9]~q  & !\prif.imemload_id [16]))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[10][9]~q ),
	.datac(\reg_file[8][9]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux54~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~12 .lut_mask = 16'hAAD8;
defparam \Mux54~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N26
cycloneive_lcell_comb \Mux36~2 (
// Equation(s):
// \Mux36~2_combout  = (\prif.imemload_id [18] & (((\reg_file[22][27]~q ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\reg_file[18][27]~q  & ((!\prif.imemload_id [19]))))

	.dataa(\reg_file[18][27]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[22][27]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux36~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~2 .lut_mask = 16'hCCE2;
defparam \Mux36~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N11
dffeas \reg_file[24][27] (
	.clk(!CLK),
	.d(\reg_file[24][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][27] .is_wysiwyg = "true";
defparam \reg_file[24][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N14
cycloneive_lcell_comb \Mux40~4 (
// Equation(s):
// \Mux40~4_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[20][23]~q ))) # (!\prif.imemload_id [18] & (\reg_file[16][23]~q ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[16][23]~q ),
	.datac(\reg_file[20][23]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux40~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~4 .lut_mask = 16'hFA44;
defparam \Mux40~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N25
dffeas \reg_file[16][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][18] .is_wysiwyg = "true";
defparam \reg_file[16][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N24
cycloneive_lcell_comb \Mux45~4 (
// Equation(s):
// \Mux45~4_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[24][18]~q )) # (!\prif.imemload_id [19] & ((\reg_file[16][18]~q )))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[24][18]~q ),
	.datac(\reg_file[16][18]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux45~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~4 .lut_mask = 16'hEE50;
defparam \Mux45~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N14
cycloneive_lcell_comb \Mux45~12 (
// Equation(s):
// \Mux45~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][18]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][18]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][18]~q ),
	.datad(\reg_file[5][18]~q ),
	.cin(gnd),
	.combout(\Mux45~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~12 .lut_mask = 16'hBA98;
defparam \Mux45~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N7
dffeas \reg_file[2][18] (
	.clk(!CLK),
	.d(\reg_file[2][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][18] .is_wysiwyg = "true";
defparam \reg_file[2][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N3
dffeas \reg_file[18][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][24] .is_wysiwyg = "true";
defparam \reg_file[18][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N31
dffeas \reg_file[20][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][24] .is_wysiwyg = "true";
defparam \reg_file[20][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N26
cycloneive_lcell_comb \Mux47~2 (
// Equation(s):
// \Mux47~2_combout  = (\prif.imemload_id [19] & (((\reg_file[26][16]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[18][16]~q  & ((!\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[18][16]~q ),
	.datac(\reg_file[26][16]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux47~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~2 .lut_mask = 16'hAAE4;
defparam \Mux47~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N17
dffeas \reg_file[26][19] (
	.clk(!CLK),
	.d(\reg_file[26][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][19] .is_wysiwyg = "true";
defparam \reg_file[26][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N1
dffeas \reg_file[20][17] (
	.clk(!CLK),
	.d(\reg_file[20][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][17] .is_wysiwyg = "true";
defparam \reg_file[20][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N6
cycloneive_lcell_comb \Mux46~4 (
// Equation(s):
// \Mux46~4_combout  = (\prif.imemload_id [18] & ((\reg_file[20][17]~q ) # ((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (((\reg_file[16][17]~q  & !\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[20][17]~q ),
	.datac(\reg_file[16][17]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux46~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~4 .lut_mask = 16'hAAD8;
defparam \Mux46~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N4
cycloneive_lcell_comb \Mux43~2 (
// Equation(s):
// \Mux43~2_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[26][20]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & ((\reg_file[18][20]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[26][20]~q ),
	.datad(\reg_file[18][20]~q ),
	.cin(gnd),
	.combout(\Mux43~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~2 .lut_mask = 16'hB9A8;
defparam \Mux43~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N31
dffeas \reg_file[8][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][20] .is_wysiwyg = "true";
defparam \reg_file[8][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N7
dffeas \reg_file[18][28] (
	.clk(!CLK),
	.d(\reg_file[18][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][28] .is_wysiwyg = "true";
defparam \reg_file[18][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N8
cycloneive_lcell_comb \Mux35~2 (
// Equation(s):
// \Mux35~2_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[26][28]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & ((\reg_file[18][28]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[26][28]~q ),
	.datad(\reg_file[18][28]~q ),
	.cin(gnd),
	.combout(\Mux35~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~2 .lut_mask = 16'hB9A8;
defparam \Mux35~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N12
cycloneive_lcell_comb \Mux35~12 (
// Equation(s):
// \Mux35~12_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & (\reg_file[5][28]~q )) # (!\prif.imemload_id [16] & ((\reg_file[4][28]~q )))))

	.dataa(\reg_file[5][28]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][28]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux35~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~12 .lut_mask = 16'hEE30;
defparam \Mux35~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N20
cycloneive_lcell_comb \Mux37~2 (
// Equation(s):
// \Mux37~2_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[26][26]~q )) # (!\prif.imemload_id [19] & ((\reg_file[18][26]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[26][26]~q ),
	.datad(\reg_file[18][26]~q ),
	.cin(gnd),
	.combout(\Mux37~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~2 .lut_mask = 16'hD9C8;
defparam \Mux37~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N7
dffeas \reg_file[24][26] (
	.clk(!CLK),
	.d(\reg_file[24][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][26] .is_wysiwyg = "true";
defparam \reg_file[24][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N10
cycloneive_lcell_comb \Mux37~4 (
// Equation(s):
// \Mux37~4_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[24][26]~q ))) # (!\prif.imemload_id [19] & (\reg_file[16][26]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[16][26]~q ),
	.datad(\reg_file[24][26]~q ),
	.cin(gnd),
	.combout(\Mux37~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~4 .lut_mask = 16'hDC98;
defparam \Mux37~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N12
cycloneive_lcell_comb \Mux38~4 (
// Equation(s):
// \Mux38~4_combout  = (\prif.imemload_id [18] & (((\reg_file[20][25]~q ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\reg_file[16][25]~q  & ((!\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[16][25]~q ),
	.datac(\reg_file[20][25]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux38~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~4 .lut_mask = 16'hAAE4;
defparam \Mux38~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N2
cycloneive_lcell_comb \Mux38~14 (
// Equation(s):
// \Mux38~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][25]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][25]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[1][25]~q ),
	.datad(\reg_file[3][25]~q ),
	.cin(gnd),
	.combout(\Mux38~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~14 .lut_mask = 16'hA820;
defparam \Mux38~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N30
cycloneive_lcell_comb \Mux29~4 (
// Equation(s):
// \Mux29~4_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[20][2]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[16][2]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][2]~q ),
	.datad(\reg_file[20][2]~q ),
	.cin(gnd),
	.combout(\Mux29~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~4 .lut_mask = 16'hBA98;
defparam \Mux29~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N26
cycloneive_lcell_comb \Mux29~12 (
// Equation(s):
// \Mux29~12_combout  = (\prif.imemload_id [22] & ((\reg_file[10][2]~q ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\reg_file[8][2]~q  & !\prif.imemload_id [21]))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[10][2]~q ),
	.datac(\reg_file[8][2]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux29~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~12 .lut_mask = 16'hAAD8;
defparam \Mux29~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N6
cycloneive_lcell_comb \Mux29~14 (
// Equation(s):
// \Mux29~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][2]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][2]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[1][2]~q ),
	.datad(\reg_file[3][2]~q ),
	.cin(gnd),
	.combout(\Mux29~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~14 .lut_mask = 16'hA820;
defparam \Mux29~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N8
cycloneive_lcell_comb \Mux27~2 (
// Equation(s):
// \Mux27~2_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\reg_file[22][4]~q )) # (!\prif.imemload_id [23] & ((\reg_file[18][4]~q )))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[22][4]~q ),
	.datac(\reg_file[18][4]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux27~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~2 .lut_mask = 16'hEE50;
defparam \Mux27~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N30
cycloneive_lcell_comb \Mux27~12 (
// Equation(s):
// \Mux27~12_combout  = (\prif.imemload_id [22] & ((\prif.imemload_id [21]) # ((\reg_file[10][4]~q )))) # (!\prif.imemload_id [22] & (!\prif.imemload_id [21] & (\reg_file[8][4]~q )))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[8][4]~q ),
	.datad(\reg_file[10][4]~q ),
	.cin(gnd),
	.combout(\Mux27~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~12 .lut_mask = 16'hBA98;
defparam \Mux27~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N12
cycloneive_lcell_comb \Mux28~14 (
// Equation(s):
// \Mux28~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][3]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][3]~q ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[1][3]~q ),
	.datac(\reg_file[3][3]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux28~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~14 .lut_mask = 16'hA088;
defparam \Mux28~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N20
cycloneive_lcell_comb \Mux23~14 (
// Equation(s):
// \Mux23~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][8]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][8]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[1][8]~q ),
	.datad(\reg_file[3][8]~q ),
	.cin(gnd),
	.combout(\Mux23~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~14 .lut_mask = 16'hA820;
defparam \Mux23~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N6
cycloneive_lcell_comb \Mux25~2 (
// Equation(s):
// \Mux25~2_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[22][6]~q ))) # (!\prif.imemload_id [23] & (\reg_file[18][6]~q ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[18][6]~q ),
	.datac(\reg_file[22][6]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux25~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~2 .lut_mask = 16'hFA44;
defparam \Mux25~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N18
cycloneive_lcell_comb \Mux15~12 (
// Equation(s):
// \Mux15~12_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[10][16]~q ))) # (!\prif.imemload_id [22] & (\reg_file[8][16]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[8][16]~q ),
	.datad(\reg_file[10][16]~q ),
	.cin(gnd),
	.combout(\Mux15~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~12 .lut_mask = 16'hDC98;
defparam \Mux15~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N20
cycloneive_lcell_comb \Mux17~14 (
// Equation(s):
// \Mux17~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][14]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][14]~q ))))

	.dataa(\reg_file[1][14]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][14]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux17~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~14 .lut_mask = 16'hE200;
defparam \Mux17~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N8
cycloneive_lcell_comb \Mux18~12 (
// Equation(s):
// \Mux18~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][13]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[4][13]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[4][13]~q ),
	.datad(\reg_file[5][13]~q ),
	.cin(gnd),
	.combout(\Mux18~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~12 .lut_mask = 16'hBA98;
defparam \Mux18~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N22
cycloneive_lcell_comb \Mux19~2 (
// Equation(s):
// \Mux19~2_combout  = (\prif.imemload_id [23] & (((\reg_file[22][12]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[18][12]~q  & ((!\prif.imemload_id [24]))))

	.dataa(\reg_file[18][12]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[22][12]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux19~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~2 .lut_mask = 16'hCCE2;
defparam \Mux19~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N14
cycloneive_lcell_comb \Mux19~12 (
// Equation(s):
// \Mux19~12_combout  = (\prif.imemload_id [22] & ((\reg_file[10][12]~q ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\reg_file[8][12]~q  & !\prif.imemload_id [21]))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[10][12]~q ),
	.datac(\reg_file[8][12]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux19~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~12 .lut_mask = 16'hAAD8;
defparam \Mux19~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N2
cycloneive_lcell_comb \Mux19~14 (
// Equation(s):
// \Mux19~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][12]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][12]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][12]~q ),
	.datad(\reg_file[1][12]~q ),
	.cin(gnd),
	.combout(\Mux19~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~14 .lut_mask = 16'hA280;
defparam \Mux19~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N2
cycloneive_lcell_comb \Mux21~12 (
// Equation(s):
// \Mux21~12_combout  = (\prif.imemload_id [22] & ((\prif.imemload_id [21]) # ((\reg_file[10][10]~q )))) # (!\prif.imemload_id [22] & (!\prif.imemload_id [21] & (\reg_file[8][10]~q )))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[8][10]~q ),
	.datad(\reg_file[10][10]~q ),
	.cin(gnd),
	.combout(\Mux21~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~12 .lut_mask = 16'hBA98;
defparam \Mux21~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N0
cycloneive_lcell_comb \Mux22~2 (
// Equation(s):
// \Mux22~2_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[26][9]~q ))) # (!\prif.imemload_id [24] & (\reg_file[18][9]~q ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[18][9]~q ),
	.datac(\reg_file[26][9]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux22~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~2 .lut_mask = 16'hFA44;
defparam \Mux22~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N14
cycloneive_lcell_comb \Mux22~14 (
// Equation(s):
// \Mux22~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][9]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][9]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[1][9]~q ),
	.datad(\reg_file[3][9]~q ),
	.cin(gnd),
	.combout(\Mux22~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~14 .lut_mask = 16'hA820;
defparam \Mux22~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N22
cycloneive_lcell_comb \Mux13~4 (
// Equation(s):
// \Mux13~4_combout  = (\prif.imemload_id [23] & (((\reg_file[20][18]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[16][18]~q  & ((!\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[16][18]~q ),
	.datac(\reg_file[20][18]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux13~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~4 .lut_mask = 16'hAAE4;
defparam \Mux13~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N18
cycloneive_lcell_comb \Mux13~12 (
// Equation(s):
// \Mux13~12_combout  = (\prif.imemload_id [22] & ((\prif.imemload_id [21]) # ((\reg_file[10][18]~q )))) # (!\prif.imemload_id [22] & (!\prif.imemload_id [21] & (\reg_file[8][18]~q )))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[8][18]~q ),
	.datad(\reg_file[10][18]~q ),
	.cin(gnd),
	.combout(\Mux13~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~12 .lut_mask = 16'hBA98;
defparam \Mux13~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N2
cycloneive_lcell_comb \Mux14~12 (
// Equation(s):
// \Mux14~12_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[5][17]~q ))) # (!\prif.imemload_id [21] & (\reg_file[4][17]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[4][17]~q ),
	.datad(\reg_file[5][17]~q ),
	.cin(gnd),
	.combout(\Mux14~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~12 .lut_mask = 16'hDC98;
defparam \Mux14~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N26
cycloneive_lcell_comb \Mux14~14 (
// Equation(s):
// \Mux14~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][17]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][17]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[1][17]~q ),
	.datad(\reg_file[3][17]~q ),
	.cin(gnd),
	.combout(\Mux14~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~14 .lut_mask = 16'hA820;
defparam \Mux14~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N30
cycloneive_lcell_comb \Mux11~12 (
// Equation(s):
// \Mux11~12_combout  = (\prif.imemload_id [22] & ((\reg_file[10][20]~q ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\reg_file[8][20]~q  & !\prif.imemload_id [21]))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[10][20]~q ),
	.datac(\reg_file[8][20]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux11~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~12 .lut_mask = 16'hAAD8;
defparam \Mux11~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N14
cycloneive_lcell_comb \Mux11~14 (
// Equation(s):
// \Mux11~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][20]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][20]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][20]~q ),
	.datad(\reg_file[1][20]~q ),
	.cin(gnd),
	.combout(\Mux11~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~14 .lut_mask = 16'hA280;
defparam \Mux11~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N22
cycloneive_lcell_comb \Mux12~2 (
// Equation(s):
// \Mux12~2_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[26][19]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[18][19]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[18][19]~q ),
	.datad(\reg_file[26][19]~q ),
	.cin(gnd),
	.combout(\Mux12~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~2 .lut_mask = 16'hBA98;
defparam \Mux12~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N2
cycloneive_lcell_comb \Mux7~2 (
// Equation(s):
// \Mux7~2_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[22][24]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[18][24]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[18][24]~q ),
	.datad(\reg_file[22][24]~q ),
	.cin(gnd),
	.combout(\Mux7~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~2 .lut_mask = 16'hBA98;
defparam \Mux7~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N30
cycloneive_lcell_comb \Mux7~4 (
// Equation(s):
// \Mux7~4_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[20][24]~q ))) # (!\prif.imemload_id [23] & (\reg_file[16][24]~q ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[16][24]~q ),
	.datac(\reg_file[20][24]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux7~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~4 .lut_mask = 16'hFA44;
defparam \Mux7~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N8
cycloneive_lcell_comb \Mux7~12 (
// Equation(s):
// \Mux7~12_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[10][24]~q )) # (!\prif.imemload_id [22] & ((\reg_file[8][24]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[10][24]~q ),
	.datad(\reg_file[8][24]~q ),
	.cin(gnd),
	.combout(\Mux7~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~12 .lut_mask = 16'hD9C8;
defparam \Mux7~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N12
cycloneive_lcell_comb \Mux7~14 (
// Equation(s):
// \Mux7~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][24]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][24]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[1][24]~q ),
	.datad(\reg_file[3][24]~q ),
	.cin(gnd),
	.combout(\Mux7~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~14 .lut_mask = 16'hC840;
defparam \Mux7~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N18
cycloneive_lcell_comb \Mux0~2 (
// Equation(s):
// \Mux0~2_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[26][31]~q )) # (!\prif.imemload_id [24] & ((\reg_file[18][31]~q )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[26][31]~q ),
	.datad(\reg_file[18][31]~q ),
	.cin(gnd),
	.combout(\Mux0~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~2 .lut_mask = 16'hD9C8;
defparam \Mux0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N24
cycloneive_lcell_comb \Mux1~2 (
// Equation(s):
// \Mux1~2_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[22][30]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & ((\reg_file[18][30]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[22][30]~q ),
	.datad(\reg_file[18][30]~q ),
	.cin(gnd),
	.combout(\Mux1~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~2 .lut_mask = 16'hB9A8;
defparam \Mux1~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N14
cycloneive_lcell_comb \Mux1~12 (
// Equation(s):
// \Mux1~12_combout  = (\prif.imemload_id [22] & ((\reg_file[10][30]~q ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\reg_file[8][30]~q  & !\prif.imemload_id [21]))))

	.dataa(\reg_file[10][30]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[8][30]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux1~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~12 .lut_mask = 16'hCCB8;
defparam \Mux1~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N20
cycloneive_lcell_comb \Mux2~2 (
// Equation(s):
// \Mux2~2_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[26][29]~q )) # (!\prif.imemload_id [24] & ((\reg_file[18][29]~q )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[26][29]~q ),
	.datad(\reg_file[18][29]~q ),
	.cin(gnd),
	.combout(\Mux2~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~2 .lut_mask = 16'hD9C8;
defparam \Mux2~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N22
cycloneive_lcell_comb \Mux6~2 (
// Equation(s):
// \Mux6~2_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23]) # (\reg_file[26][25]~q )))) # (!\prif.imemload_id [24] & (\reg_file[18][25]~q  & (!\prif.imemload_id [23])))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[18][25]~q ),
	.datac(prifimemload_id_23),
	.datad(\reg_file[26][25]~q ),
	.cin(gnd),
	.combout(\Mux6~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~2 .lut_mask = 16'hAEA4;
defparam \Mux6~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N4
cycloneive_lcell_comb \Mux3~2 (
// Equation(s):
// \Mux3~2_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[22][28]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[18][28]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[18][28]~q ),
	.datad(\reg_file[22][28]~q ),
	.cin(gnd),
	.combout(\Mux3~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~2 .lut_mask = 16'hBA98;
defparam \Mux3~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N10
cycloneive_lcell_comb \Mux3~4 (
// Equation(s):
// \Mux3~4_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[20][28]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & ((\reg_file[16][28]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[20][28]~q ),
	.datad(\reg_file[16][28]~q ),
	.cin(gnd),
	.combout(\Mux3~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~4 .lut_mask = 16'hB9A8;
defparam \Mux3~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N10
cycloneive_lcell_comb \reg_file[24][27]~feeder (
// Equation(s):
// \reg_file[24][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][27]~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[24][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][27]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[24][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N6
cycloneive_lcell_comb \reg_file[2][18]~feeder (
// Equation(s):
// \reg_file[2][18]~feeder_combout  = \reg_file_nxt[31][18]~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][18]~83_combout ),
	.cin(gnd),
	.combout(\reg_file[2][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][18]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[2][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N16
cycloneive_lcell_comb \reg_file[26][19]~feeder (
// Equation(s):
// \reg_file[26][19]~feeder_combout  = \reg_file_nxt[31][19]~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][19]~86_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[26][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[26][19]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[26][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N0
cycloneive_lcell_comb \reg_file[20][17]~feeder (
// Equation(s):
// \reg_file[20][17]~feeder_combout  = \reg_file_nxt[31][17]~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][17]~87_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[20][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[20][17]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[20][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N6
cycloneive_lcell_comb \reg_file[18][28]~feeder (
// Equation(s):
// \reg_file[18][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][28]~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[18][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[18][28]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[18][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N6
cycloneive_lcell_comb \reg_file[24][26]~feeder (
// Equation(s):
// \reg_file[24][26]~feeder_combout  = \reg_file_nxt[31][26]~91_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][26]~91_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[24][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][26]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[24][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N14
cycloneive_lcell_comb \Mux62~9 (
// Equation(s):
// Mux62 = (\prif.imemload_id [16] & ((\Mux62~6_combout  & ((\Mux62~8_combout ))) # (!\Mux62~6_combout  & (\Mux62~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux62~6_combout ))))

	.dataa(\Mux62~1_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux62~6_combout ),
	.datad(\Mux62~8_combout ),
	.cin(gnd),
	.combout(Mux62),
	.cout());
// synopsys translate_off
defparam \Mux62~9 .lut_mask = 16'hF838;
defparam \Mux62~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N12
cycloneive_lcell_comb \Mux62~19 (
// Equation(s):
// Mux621 = (\Mux62~16_combout  & ((\Mux62~18_combout ) # ((!\prif.imemload_id [18])))) # (!\Mux62~16_combout  & (((\prif.imemload_id [18] & \Mux62~11_combout ))))

	.dataa(\Mux62~16_combout ),
	.datab(\Mux62~18_combout ),
	.datac(prifimemload_id_18),
	.datad(\Mux62~11_combout ),
	.cin(gnd),
	.combout(Mux621),
	.cout());
// synopsys translate_off
defparam \Mux62~19 .lut_mask = 16'hDA8A;
defparam \Mux62~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N8
cycloneive_lcell_comb \Mux30~9 (
// Equation(s):
// Mux30 = (\prif.imemload_id [21] & ((\Mux30~6_combout  & ((\Mux30~8_combout ))) # (!\Mux30~6_combout  & (\Mux30~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux30~6_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\Mux30~1_combout ),
	.datac(\Mux30~8_combout ),
	.datad(\Mux30~6_combout ),
	.cin(gnd),
	.combout(Mux30),
	.cout());
// synopsys translate_off
defparam \Mux30~9 .lut_mask = 16'hF588;
defparam \Mux30~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N22
cycloneive_lcell_comb \Mux30~19 (
// Equation(s):
// Mux301 = (\Mux30~16_combout  & (((\Mux30~18_combout )) # (!\prif.imemload_id [24]))) # (!\Mux30~16_combout  & (\prif.imemload_id [24] & (\Mux30~11_combout )))

	.dataa(\Mux30~16_combout ),
	.datab(prifimemload_id_24),
	.datac(\Mux30~11_combout ),
	.datad(\Mux30~18_combout ),
	.cin(gnd),
	.combout(Mux301),
	.cout());
// synopsys translate_off
defparam \Mux30~19 .lut_mask = 16'hEA62;
defparam \Mux30~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N20
cycloneive_lcell_comb \Mux63~9 (
// Equation(s):
// Mux63 = (\prif.imemload_id [16] & ((\Mux63~6_combout  & (\Mux63~8_combout )) # (!\Mux63~6_combout  & ((\Mux63~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux63~6_combout ))))

	.dataa(\Mux63~8_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux63~1_combout ),
	.datad(\Mux63~6_combout ),
	.cin(gnd),
	.combout(Mux63),
	.cout());
// synopsys translate_off
defparam \Mux63~9 .lut_mask = 16'hBBC0;
defparam \Mux63~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N30
cycloneive_lcell_comb \Mux63~19 (
// Equation(s):
// Mux631 = (\Mux63~16_combout  & ((\Mux63~18_combout ) # ((!\prif.imemload_id [19])))) # (!\Mux63~16_combout  & (((\Mux63~11_combout  & \prif.imemload_id [19]))))

	.dataa(\Mux63~18_combout ),
	.datab(\Mux63~16_combout ),
	.datac(\Mux63~11_combout ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(Mux631),
	.cout());
// synopsys translate_off
defparam \Mux63~19 .lut_mask = 16'hB8CC;
defparam \Mux63~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N6
cycloneive_lcell_comb \Mux31~9 (
// Equation(s):
// Mux31 = (\Mux31~6_combout  & ((\Mux31~8_combout ) # ((!\prif.imemload_id [21])))) # (!\Mux31~6_combout  & (((\prif.imemload_id [21] & \Mux31~1_combout ))))

	.dataa(\Mux31~8_combout ),
	.datab(\Mux31~6_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux31~1_combout ),
	.cin(gnd),
	.combout(Mux31),
	.cout());
// synopsys translate_off
defparam \Mux31~9 .lut_mask = 16'hBC8C;
defparam \Mux31~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N4
cycloneive_lcell_comb \Mux31~19 (
// Equation(s):
// Mux311 = (\prif.imemload_id [23] & ((\Mux31~16_combout  & (\Mux31~18_combout )) # (!\Mux31~16_combout  & ((\Mux31~11_combout ))))) # (!\prif.imemload_id [23] & (\Mux31~16_combout ))

	.dataa(prifimemload_id_23),
	.datab(\Mux31~16_combout ),
	.datac(\Mux31~18_combout ),
	.datad(\Mux31~11_combout ),
	.cin(gnd),
	.combout(Mux311),
	.cout());
// synopsys translate_off
defparam \Mux31~19 .lut_mask = 16'hE6C4;
defparam \Mux31~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N2
cycloneive_lcell_comb \Mux60~9 (
// Equation(s):
// Mux60 = (\prif.imemload_id [16] & ((\Mux60~6_combout  & (\Mux60~8_combout )) # (!\Mux60~6_combout  & ((\Mux60~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux60~6_combout ))))

	.dataa(\Mux60~8_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux60~1_combout ),
	.datad(\Mux60~6_combout ),
	.cin(gnd),
	.combout(Mux60),
	.cout());
// synopsys translate_off
defparam \Mux60~9 .lut_mask = 16'hBBC0;
defparam \Mux60~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N4
cycloneive_lcell_comb \Mux60~19 (
// Equation(s):
// Mux601 = (\prif.imemload_id [18] & ((\Mux60~16_combout  & (\Mux60~18_combout )) # (!\Mux60~16_combout  & ((\Mux60~11_combout ))))) # (!\prif.imemload_id [18] & (((\Mux60~16_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux60~18_combout ),
	.datac(\Mux60~16_combout ),
	.datad(\Mux60~11_combout ),
	.cin(gnd),
	.combout(Mux601),
	.cout());
// synopsys translate_off
defparam \Mux60~19 .lut_mask = 16'hDAD0;
defparam \Mux60~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N24
cycloneive_lcell_comb \Mux61~9 (
// Equation(s):
// Mux61 = (\Mux61~6_combout  & ((\Mux61~8_combout ) # ((!\prif.imemload_id [16])))) # (!\Mux61~6_combout  & (((\prif.imemload_id [16] & \Mux61~1_combout ))))

	.dataa(\Mux61~6_combout ),
	.datab(\Mux61~8_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux61~1_combout ),
	.cin(gnd),
	.combout(Mux61),
	.cout());
// synopsys translate_off
defparam \Mux61~9 .lut_mask = 16'hDA8A;
defparam \Mux61~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N18
cycloneive_lcell_comb \Mux61~19 (
// Equation(s):
// Mux611 = (\prif.imemload_id [19] & ((\Mux61~16_combout  & ((\Mux61~18_combout ))) # (!\Mux61~16_combout  & (\Mux61~11_combout )))) # (!\prif.imemload_id [19] & (((\Mux61~16_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\Mux61~11_combout ),
	.datac(\Mux61~18_combout ),
	.datad(\Mux61~16_combout ),
	.cin(gnd),
	.combout(Mux611),
	.cout());
// synopsys translate_off
defparam \Mux61~19 .lut_mask = 16'hF588;
defparam \Mux61~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N26
cycloneive_lcell_comb \Mux59~9 (
// Equation(s):
// Mux59 = (\Mux59~6_combout  & ((\Mux59~8_combout ) # ((!\prif.imemload_id [16])))) # (!\Mux59~6_combout  & (((\prif.imemload_id [16] & \Mux59~1_combout ))))

	.dataa(\Mux59~8_combout ),
	.datab(\Mux59~6_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux59~1_combout ),
	.cin(gnd),
	.combout(Mux59),
	.cout());
// synopsys translate_off
defparam \Mux59~9 .lut_mask = 16'hBC8C;
defparam \Mux59~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N0
cycloneive_lcell_comb \Mux59~19 (
// Equation(s):
// Mux591 = (\prif.imemload_id [19] & ((\Mux59~16_combout  & ((\Mux59~18_combout ))) # (!\Mux59~16_combout  & (\Mux59~11_combout )))) # (!\prif.imemload_id [19] & (((\Mux59~16_combout ))))

	.dataa(\Mux59~11_combout ),
	.datab(prifimemload_id_19),
	.datac(\Mux59~16_combout ),
	.datad(\Mux59~18_combout ),
	.cin(gnd),
	.combout(Mux591),
	.cout());
// synopsys translate_off
defparam \Mux59~19 .lut_mask = 16'hF838;
defparam \Mux59~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N16
cycloneive_lcell_comb \Mux32~9 (
// Equation(s):
// Mux32 = (\prif.imemload_id [16] & ((\Mux32~6_combout  & ((\Mux32~8_combout ))) # (!\Mux32~6_combout  & (\Mux32~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux32~6_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\Mux32~1_combout ),
	.datac(\Mux32~6_combout ),
	.datad(\Mux32~8_combout ),
	.cin(gnd),
	.combout(Mux32),
	.cout());
// synopsys translate_off
defparam \Mux32~9 .lut_mask = 16'hF858;
defparam \Mux32~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N8
cycloneive_lcell_comb \Mux32~19 (
// Equation(s):
// Mux321 = (\prif.imemload_id [18] & ((\Mux32~16_combout  & (\Mux32~18_combout )) # (!\Mux32~16_combout  & ((\Mux32~11_combout ))))) # (!\prif.imemload_id [18] & (((\Mux32~16_combout ))))

	.dataa(\Mux32~18_combout ),
	.datab(\Mux32~11_combout ),
	.datac(prifimemload_id_18),
	.datad(\Mux32~16_combout ),
	.cin(gnd),
	.combout(Mux321),
	.cout());
// synopsys translate_off
defparam \Mux32~19 .lut_mask = 16'hAFC0;
defparam \Mux32~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N22
cycloneive_lcell_comb \Mux33~9 (
// Equation(s):
// Mux33 = (\prif.imemload_id [16] & ((\Mux33~6_combout  & (\Mux33~8_combout )) # (!\Mux33~6_combout  & ((\Mux33~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux33~6_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\Mux33~8_combout ),
	.datac(\Mux33~1_combout ),
	.datad(\Mux33~6_combout ),
	.cin(gnd),
	.combout(Mux33),
	.cout());
// synopsys translate_off
defparam \Mux33~9 .lut_mask = 16'hDDA0;
defparam \Mux33~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N6
cycloneive_lcell_comb \Mux33~19 (
// Equation(s):
// Mux331 = (\Mux33~16_combout  & ((\Mux33~18_combout ) # ((!\prif.imemload_id [19])))) # (!\Mux33~16_combout  & (((\prif.imemload_id [19] & \Mux33~11_combout ))))

	.dataa(\Mux33~16_combout ),
	.datab(\Mux33~18_combout ),
	.datac(prifimemload_id_19),
	.datad(\Mux33~11_combout ),
	.cin(gnd),
	.combout(Mux331),
	.cout());
// synopsys translate_off
defparam \Mux33~19 .lut_mask = 16'hDA8A;
defparam \Mux33~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N2
cycloneive_lcell_comb \Mux34~9 (
// Equation(s):
// Mux34 = (\prif.imemload_id [16] & ((\Mux34~6_combout  & (\Mux34~8_combout )) # (!\Mux34~6_combout  & ((\Mux34~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux34~6_combout ))))

	.dataa(\Mux34~8_combout ),
	.datab(\Mux34~1_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux34~6_combout ),
	.cin(gnd),
	.combout(Mux34),
	.cout());
// synopsys translate_off
defparam \Mux34~9 .lut_mask = 16'hAFC0;
defparam \Mux34~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N2
cycloneive_lcell_comb \Mux34~19 (
// Equation(s):
// Mux341 = (\prif.imemload_id [18] & ((\Mux34~16_combout  & (\Mux34~18_combout )) # (!\Mux34~16_combout  & ((\Mux34~11_combout ))))) # (!\prif.imemload_id [18] & (((\Mux34~16_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux34~18_combout ),
	.datac(\Mux34~16_combout ),
	.datad(\Mux34~11_combout ),
	.cin(gnd),
	.combout(Mux341),
	.cout());
// synopsys translate_off
defparam \Mux34~19 .lut_mask = 16'hDAD0;
defparam \Mux34~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N16
cycloneive_lcell_comb \Mux58~9 (
// Equation(s):
// Mux58 = (\prif.imemload_id [16] & ((\Mux58~6_combout  & ((\Mux58~8_combout ))) # (!\Mux58~6_combout  & (\Mux58~1_combout )))) # (!\prif.imemload_id [16] & (\Mux58~6_combout ))

	.dataa(prifimemload_id_16),
	.datab(\Mux58~6_combout ),
	.datac(\Mux58~1_combout ),
	.datad(\Mux58~8_combout ),
	.cin(gnd),
	.combout(Mux58),
	.cout());
// synopsys translate_off
defparam \Mux58~9 .lut_mask = 16'hEC64;
defparam \Mux58~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N24
cycloneive_lcell_comb \Mux58~19 (
// Equation(s):
// Mux581 = (\prif.imemload_id [18] & ((\Mux58~16_combout  & ((\Mux58~18_combout ))) # (!\Mux58~16_combout  & (\Mux58~11_combout )))) # (!\prif.imemload_id [18] & (((\Mux58~16_combout ))))

	.dataa(\Mux58~11_combout ),
	.datab(prifimemload_id_18),
	.datac(\Mux58~16_combout ),
	.datad(\Mux58~18_combout ),
	.cin(gnd),
	.combout(Mux581),
	.cout());
// synopsys translate_off
defparam \Mux58~19 .lut_mask = 16'hF838;
defparam \Mux58~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N8
cycloneive_lcell_comb \Mux48~9 (
// Equation(s):
// Mux48 = (\prif.imemload_id [16] & ((\Mux48~6_combout  & ((\Mux48~8_combout ))) # (!\Mux48~6_combout  & (\Mux48~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux48~6_combout ))))

	.dataa(\Mux48~1_combout ),
	.datab(\Mux48~8_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux48~6_combout ),
	.cin(gnd),
	.combout(Mux48),
	.cout());
// synopsys translate_off
defparam \Mux48~9 .lut_mask = 16'hCFA0;
defparam \Mux48~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N16
cycloneive_lcell_comb \Mux48~19 (
// Equation(s):
// Mux481 = (\Mux48~16_combout  & (((\Mux48~18_combout ) # (!\prif.imemload_id [18])))) # (!\Mux48~16_combout  & (\Mux48~11_combout  & ((\prif.imemload_id [18]))))

	.dataa(\Mux48~16_combout ),
	.datab(\Mux48~11_combout ),
	.datac(\Mux48~18_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(Mux481),
	.cout());
// synopsys translate_off
defparam \Mux48~19 .lut_mask = 16'hE4AA;
defparam \Mux48~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N28
cycloneive_lcell_comb \Mux49~9 (
// Equation(s):
// Mux49 = (\Mux49~6_combout  & (((\Mux49~8_combout )) # (!\prif.imemload_id [16]))) # (!\Mux49~6_combout  & (\prif.imemload_id [16] & ((\Mux49~1_combout ))))

	.dataa(\Mux49~6_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux49~8_combout ),
	.datad(\Mux49~1_combout ),
	.cin(gnd),
	.combout(Mux49),
	.cout());
// synopsys translate_off
defparam \Mux49~9 .lut_mask = 16'hE6A2;
defparam \Mux49~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N12
cycloneive_lcell_comb \Mux49~19 (
// Equation(s):
// Mux491 = (\Mux49~16_combout  & ((\Mux49~18_combout ) # ((!\prif.imemload_id [19])))) # (!\Mux49~16_combout  & (((\Mux49~11_combout  & \prif.imemload_id [19]))))

	.dataa(\Mux49~18_combout ),
	.datab(\Mux49~11_combout ),
	.datac(\Mux49~16_combout ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(Mux491),
	.cout());
// synopsys translate_off
defparam \Mux49~19 .lut_mask = 16'hACF0;
defparam \Mux49~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N0
cycloneive_lcell_comb \Mux50~9 (
// Equation(s):
// Mux50 = (\Mux50~6_combout  & (((\Mux50~8_combout )) # (!\prif.imemload_id [16]))) # (!\Mux50~6_combout  & (\prif.imemload_id [16] & (\Mux50~1_combout )))

	.dataa(\Mux50~6_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux50~1_combout ),
	.datad(\Mux50~8_combout ),
	.cin(gnd),
	.combout(Mux50),
	.cout());
// synopsys translate_off
defparam \Mux50~9 .lut_mask = 16'hEA62;
defparam \Mux50~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N26
cycloneive_lcell_comb \Mux50~19 (
// Equation(s):
// Mux501 = (\prif.imemload_id [18] & ((\Mux50~16_combout  & ((\Mux50~18_combout ))) # (!\Mux50~16_combout  & (\Mux50~11_combout )))) # (!\prif.imemload_id [18] & (((\Mux50~16_combout ))))

	.dataa(\Mux50~11_combout ),
	.datab(\Mux50~18_combout ),
	.datac(prifimemload_id_18),
	.datad(\Mux50~16_combout ),
	.cin(gnd),
	.combout(Mux501),
	.cout());
// synopsys translate_off
defparam \Mux50~19 .lut_mask = 16'hCFA0;
defparam \Mux50~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y28_N16
cycloneive_lcell_comb \Mux51~9 (
// Equation(s):
// Mux51 = (\prif.imemload_id [16] & ((\Mux51~6_combout  & (\Mux51~8_combout )) # (!\Mux51~6_combout  & ((\Mux51~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux51~6_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\Mux51~8_combout ),
	.datac(\Mux51~6_combout ),
	.datad(\Mux51~1_combout ),
	.cin(gnd),
	.combout(Mux51),
	.cout());
// synopsys translate_off
defparam \Mux51~9 .lut_mask = 16'hDAD0;
defparam \Mux51~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N30
cycloneive_lcell_comb \Mux51~19 (
// Equation(s):
// Mux511 = (\Mux51~16_combout  & (((\Mux51~18_combout ) # (!\prif.imemload_id [19])))) # (!\Mux51~16_combout  & (\Mux51~11_combout  & ((\prif.imemload_id [19]))))

	.dataa(\Mux51~11_combout ),
	.datab(\Mux51~16_combout ),
	.datac(\Mux51~18_combout ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(Mux511),
	.cout());
// synopsys translate_off
defparam \Mux51~19 .lut_mask = 16'hE2CC;
defparam \Mux51~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N0
cycloneive_lcell_comb \Mux52~9 (
// Equation(s):
// Mux52 = (\prif.imemload_id [16] & ((\Mux52~6_combout  & (\Mux52~8_combout )) # (!\Mux52~6_combout  & ((\Mux52~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux52~6_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\Mux52~8_combout ),
	.datac(\Mux52~1_combout ),
	.datad(\Mux52~6_combout ),
	.cin(gnd),
	.combout(Mux52),
	.cout());
// synopsys translate_off
defparam \Mux52~9 .lut_mask = 16'hDDA0;
defparam \Mux52~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N22
cycloneive_lcell_comb \Mux52~19 (
// Equation(s):
// Mux521 = (\prif.imemload_id [18] & ((\Mux52~16_combout  & ((\Mux52~18_combout ))) # (!\Mux52~16_combout  & (\Mux52~11_combout )))) # (!\prif.imemload_id [18] & (\Mux52~16_combout ))

	.dataa(prifimemload_id_18),
	.datab(\Mux52~16_combout ),
	.datac(\Mux52~11_combout ),
	.datad(\Mux52~18_combout ),
	.cin(gnd),
	.combout(Mux521),
	.cout());
// synopsys translate_off
defparam \Mux52~19 .lut_mask = 16'hEC64;
defparam \Mux52~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N12
cycloneive_lcell_comb \Mux53~9 (
// Equation(s):
// Mux53 = (\prif.imemload_id [16] & ((\Mux53~6_combout  & ((\Mux53~8_combout ))) # (!\Mux53~6_combout  & (\Mux53~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux53~6_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\Mux53~1_combout ),
	.datac(\Mux53~6_combout ),
	.datad(\Mux53~8_combout ),
	.cin(gnd),
	.combout(Mux53),
	.cout());
// synopsys translate_off
defparam \Mux53~9 .lut_mask = 16'hF858;
defparam \Mux53~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N14
cycloneive_lcell_comb \Mux53~19 (
// Equation(s):
// Mux531 = (\prif.imemload_id [19] & ((\Mux53~16_combout  & (\Mux53~18_combout )) # (!\Mux53~16_combout  & ((\Mux53~11_combout ))))) # (!\prif.imemload_id [19] & (((\Mux53~16_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\Mux53~18_combout ),
	.datac(\Mux53~11_combout ),
	.datad(\Mux53~16_combout ),
	.cin(gnd),
	.combout(Mux531),
	.cout());
// synopsys translate_off
defparam \Mux53~19 .lut_mask = 16'hDDA0;
defparam \Mux53~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N22
cycloneive_lcell_comb \Mux54~9 (
// Equation(s):
// Mux54 = (\Mux54~6_combout  & (((\Mux54~8_combout )) # (!\prif.imemload_id [16]))) # (!\Mux54~6_combout  & (\prif.imemload_id [16] & (\Mux54~1_combout )))

	.dataa(\Mux54~6_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux54~1_combout ),
	.datad(\Mux54~8_combout ),
	.cin(gnd),
	.combout(Mux54),
	.cout());
// synopsys translate_off
defparam \Mux54~9 .lut_mask = 16'hEA62;
defparam \Mux54~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N20
cycloneive_lcell_comb \Mux54~19 (
// Equation(s):
// Mux541 = (\Mux54~16_combout  & ((\Mux54~18_combout ) # ((!\prif.imemload_id [18])))) # (!\Mux54~16_combout  & (((\Mux54~11_combout  & \prif.imemload_id [18]))))

	.dataa(\Mux54~18_combout ),
	.datab(\Mux54~16_combout ),
	.datac(\Mux54~11_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(Mux541),
	.cout());
// synopsys translate_off
defparam \Mux54~19 .lut_mask = 16'hB8CC;
defparam \Mux54~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N6
cycloneive_lcell_comb \Mux57~9 (
// Equation(s):
// Mux57 = (\prif.imemload_id [16] & ((\Mux57~6_combout  & ((\Mux57~8_combout ))) # (!\Mux57~6_combout  & (\Mux57~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux57~6_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\Mux57~1_combout ),
	.datac(\Mux57~8_combout ),
	.datad(\Mux57~6_combout ),
	.cin(gnd),
	.combout(Mux57),
	.cout());
// synopsys translate_off
defparam \Mux57~9 .lut_mask = 16'hF588;
defparam \Mux57~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N18
cycloneive_lcell_comb \Mux57~19 (
// Equation(s):
// Mux571 = (\Mux57~16_combout  & (((\Mux57~18_combout )) # (!\prif.imemload_id [19]))) # (!\Mux57~16_combout  & (\prif.imemload_id [19] & (\Mux57~11_combout )))

	.dataa(\Mux57~16_combout ),
	.datab(prifimemload_id_19),
	.datac(\Mux57~11_combout ),
	.datad(\Mux57~18_combout ),
	.cin(gnd),
	.combout(Mux571),
	.cout());
// synopsys translate_off
defparam \Mux57~19 .lut_mask = 16'hEA62;
defparam \Mux57~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N6
cycloneive_lcell_comb \Mux36~9 (
// Equation(s):
// Mux36 = (\prif.imemload_id [16] & ((\Mux36~6_combout  & ((\Mux36~8_combout ))) # (!\Mux36~6_combout  & (\Mux36~1_combout )))) # (!\prif.imemload_id [16] & (\Mux36~6_combout ))

	.dataa(prifimemload_id_16),
	.datab(\Mux36~6_combout ),
	.datac(\Mux36~1_combout ),
	.datad(\Mux36~8_combout ),
	.cin(gnd),
	.combout(Mux36),
	.cout());
// synopsys translate_off
defparam \Mux36~9 .lut_mask = 16'hEC64;
defparam \Mux36~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N4
cycloneive_lcell_comb \Mux36~19 (
// Equation(s):
// Mux361 = (\prif.imemload_id [18] & ((\Mux36~16_combout  & (\Mux36~18_combout )) # (!\Mux36~16_combout  & ((\Mux36~11_combout ))))) # (!\prif.imemload_id [18] & (((\Mux36~16_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux36~18_combout ),
	.datac(\Mux36~16_combout ),
	.datad(\Mux36~11_combout ),
	.cin(gnd),
	.combout(Mux361),
	.cout());
// synopsys translate_off
defparam \Mux36~19 .lut_mask = 16'hDAD0;
defparam \Mux36~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N30
cycloneive_lcell_comb \Mux40~9 (
// Equation(s):
// Mux40 = (\Mux40~6_combout  & (((\Mux40~8_combout ) # (!\prif.imemload_id [16])))) # (!\Mux40~6_combout  & (\Mux40~1_combout  & (\prif.imemload_id [16])))

	.dataa(\Mux40~1_combout ),
	.datab(\Mux40~6_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux40~8_combout ),
	.cin(gnd),
	.combout(Mux40),
	.cout());
// synopsys translate_off
defparam \Mux40~9 .lut_mask = 16'hEC2C;
defparam \Mux40~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N18
cycloneive_lcell_comb \Mux40~19 (
// Equation(s):
// Mux401 = (\prif.imemload_id [18] & ((\Mux40~16_combout  & (\Mux40~18_combout )) # (!\Mux40~16_combout  & ((\Mux40~11_combout ))))) # (!\prif.imemload_id [18] & (((\Mux40~16_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux40~18_combout ),
	.datac(\Mux40~11_combout ),
	.datad(\Mux40~16_combout ),
	.cin(gnd),
	.combout(Mux401),
	.cout());
// synopsys translate_off
defparam \Mux40~19 .lut_mask = 16'hDDA0;
defparam \Mux40~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N4
cycloneive_lcell_comb \Mux45~9 (
// Equation(s):
// Mux45 = (\Mux45~6_combout  & (((\Mux45~8_combout )) # (!\prif.imemload_id [16]))) # (!\Mux45~6_combout  & (\prif.imemload_id [16] & ((\Mux45~1_combout ))))

	.dataa(\Mux45~6_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux45~8_combout ),
	.datad(\Mux45~1_combout ),
	.cin(gnd),
	.combout(Mux45),
	.cout());
// synopsys translate_off
defparam \Mux45~9 .lut_mask = 16'hE6A2;
defparam \Mux45~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N28
cycloneive_lcell_comb \Mux45~19 (
// Equation(s):
// Mux451 = (\Mux45~16_combout  & (((\Mux45~18_combout )) # (!\prif.imemload_id [19]))) # (!\Mux45~16_combout  & (\prif.imemload_id [19] & ((\Mux45~11_combout ))))

	.dataa(\Mux45~16_combout ),
	.datab(prifimemload_id_19),
	.datac(\Mux45~18_combout ),
	.datad(\Mux45~11_combout ),
	.cin(gnd),
	.combout(Mux451),
	.cout());
// synopsys translate_off
defparam \Mux45~19 .lut_mask = 16'hE6A2;
defparam \Mux45~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N14
cycloneive_lcell_comb \Mux39~9 (
// Equation(s):
// Mux39 = (\prif.imemload_id [16] & ((\Mux39~6_combout  & ((\Mux39~8_combout ))) # (!\Mux39~6_combout  & (\Mux39~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux39~6_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\Mux39~1_combout ),
	.datac(\Mux39~6_combout ),
	.datad(\Mux39~8_combout ),
	.cin(gnd),
	.combout(Mux39),
	.cout());
// synopsys translate_off
defparam \Mux39~9 .lut_mask = 16'hF858;
defparam \Mux39~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N16
cycloneive_lcell_comb \Mux39~19 (
// Equation(s):
// Mux391 = (\Mux39~16_combout  & (((\Mux39~18_combout ) # (!\prif.imemload_id [19])))) # (!\Mux39~16_combout  & (\Mux39~11_combout  & (\prif.imemload_id [19])))

	.dataa(\Mux39~16_combout ),
	.datab(\Mux39~11_combout ),
	.datac(prifimemload_id_19),
	.datad(\Mux39~18_combout ),
	.cin(gnd),
	.combout(Mux391),
	.cout());
// synopsys translate_off
defparam \Mux39~19 .lut_mask = 16'hEA4A;
defparam \Mux39~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N30
cycloneive_lcell_comb \Mux47~9 (
// Equation(s):
// Mux47 = (\prif.imemload_id [16] & ((\Mux47~6_combout  & ((\Mux47~8_combout ))) # (!\Mux47~6_combout  & (\Mux47~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux47~6_combout ))))

	.dataa(\Mux47~1_combout ),
	.datab(\Mux47~8_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux47~6_combout ),
	.cin(gnd),
	.combout(Mux47),
	.cout());
// synopsys translate_off
defparam \Mux47~9 .lut_mask = 16'hCFA0;
defparam \Mux47~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N6
cycloneive_lcell_comb \Mux47~19 (
// Equation(s):
// Mux471 = (\prif.imemload_id [19] & ((\Mux47~16_combout  & (\Mux47~18_combout )) # (!\Mux47~16_combout  & ((\Mux47~11_combout ))))) # (!\prif.imemload_id [19] & (\Mux47~16_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux47~16_combout ),
	.datac(\Mux47~18_combout ),
	.datad(\Mux47~11_combout ),
	.cin(gnd),
	.combout(Mux471),
	.cout());
// synopsys translate_off
defparam \Mux47~19 .lut_mask = 16'hE6C4;
defparam \Mux47~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N12
cycloneive_lcell_comb \Mux44~9 (
// Equation(s):
// Mux44 = (\prif.imemload_id [16] & ((\Mux44~6_combout  & ((\Mux44~8_combout ))) # (!\Mux44~6_combout  & (\Mux44~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux44~6_combout ))))

	.dataa(\Mux44~1_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux44~6_combout ),
	.datad(\Mux44~8_combout ),
	.cin(gnd),
	.combout(Mux44),
	.cout());
// synopsys translate_off
defparam \Mux44~9 .lut_mask = 16'hF838;
defparam \Mux44~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N12
cycloneive_lcell_comb \Mux44~19 (
// Equation(s):
// Mux441 = (\prif.imemload_id [18] & ((\Mux44~16_combout  & ((\Mux44~18_combout ))) # (!\Mux44~16_combout  & (\Mux44~11_combout )))) # (!\prif.imemload_id [18] & (((\Mux44~16_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux44~11_combout ),
	.datac(\Mux44~18_combout ),
	.datad(\Mux44~16_combout ),
	.cin(gnd),
	.combout(Mux441),
	.cout());
// synopsys translate_off
defparam \Mux44~19 .lut_mask = 16'hF588;
defparam \Mux44~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N0
cycloneive_lcell_comb \Mux46~9 (
// Equation(s):
// Mux46 = (\prif.imemload_id [16] & ((\Mux46~6_combout  & ((\Mux46~8_combout ))) # (!\Mux46~6_combout  & (\Mux46~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux46~6_combout ))))

	.dataa(\Mux46~1_combout ),
	.datab(\Mux46~8_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux46~6_combout ),
	.cin(gnd),
	.combout(Mux46),
	.cout());
// synopsys translate_off
defparam \Mux46~9 .lut_mask = 16'hCFA0;
defparam \Mux46~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N16
cycloneive_lcell_comb \Mux46~19 (
// Equation(s):
// Mux461 = (\Mux46~16_combout  & ((\Mux46~18_combout ) # ((!\prif.imemload_id [18])))) # (!\Mux46~16_combout  & (((\Mux46~11_combout  & \prif.imemload_id [18]))))

	.dataa(\Mux46~16_combout ),
	.datab(\Mux46~18_combout ),
	.datac(\Mux46~11_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(Mux461),
	.cout());
// synopsys translate_off
defparam \Mux46~19 .lut_mask = 16'hD8AA;
defparam \Mux46~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N22
cycloneive_lcell_comb \Mux42~9 (
// Equation(s):
// Mux42 = (\prif.imemload_id [16] & ((\Mux42~6_combout  & (\Mux42~8_combout )) # (!\Mux42~6_combout  & ((\Mux42~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux42~6_combout ))))

	.dataa(\Mux42~8_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux42~1_combout ),
	.datad(\Mux42~6_combout ),
	.cin(gnd),
	.combout(Mux42),
	.cout());
// synopsys translate_off
defparam \Mux42~9 .lut_mask = 16'hBBC0;
defparam \Mux42~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N24
cycloneive_lcell_comb \Mux42~19 (
// Equation(s):
// Mux421 = (\prif.imemload_id [18] & ((\Mux42~16_combout  & (\Mux42~18_combout )) # (!\Mux42~16_combout  & ((\Mux42~11_combout ))))) # (!\prif.imemload_id [18] & (((\Mux42~16_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux42~18_combout ),
	.datac(\Mux42~11_combout ),
	.datad(\Mux42~16_combout ),
	.cin(gnd),
	.combout(Mux421),
	.cout());
// synopsys translate_off
defparam \Mux42~19 .lut_mask = 16'hDDA0;
defparam \Mux42~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N30
cycloneive_lcell_comb \Mux43~9 (
// Equation(s):
// Mux43 = (\prif.imemload_id [16] & ((\Mux43~6_combout  & (\Mux43~8_combout )) # (!\Mux43~6_combout  & ((\Mux43~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux43~6_combout ))))

	.dataa(\Mux43~8_combout ),
	.datab(\Mux43~1_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux43~6_combout ),
	.cin(gnd),
	.combout(Mux43),
	.cout());
// synopsys translate_off
defparam \Mux43~9 .lut_mask = 16'hAFC0;
defparam \Mux43~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N0
cycloneive_lcell_comb \Mux43~19 (
// Equation(s):
// Mux431 = (\prif.imemload_id [19] & ((\Mux43~16_combout  & ((\Mux43~18_combout ))) # (!\Mux43~16_combout  & (\Mux43~11_combout )))) # (!\prif.imemload_id [19] & (((\Mux43~16_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\Mux43~11_combout ),
	.datac(\Mux43~18_combout ),
	.datad(\Mux43~16_combout ),
	.cin(gnd),
	.combout(Mux431),
	.cout());
// synopsys translate_off
defparam \Mux43~19 .lut_mask = 16'hF588;
defparam \Mux43~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N8
cycloneive_lcell_comb \Mux35~9 (
// Equation(s):
// Mux35 = (\prif.imemload_id [16] & ((\Mux35~6_combout  & ((\Mux35~8_combout ))) # (!\Mux35~6_combout  & (\Mux35~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux35~6_combout ))))

	.dataa(\Mux35~1_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux35~6_combout ),
	.datad(\Mux35~8_combout ),
	.cin(gnd),
	.combout(Mux35),
	.cout());
// synopsys translate_off
defparam \Mux35~9 .lut_mask = 16'hF838;
defparam \Mux35~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N14
cycloneive_lcell_comb \Mux35~19 (
// Equation(s):
// Mux351 = (\prif.imemload_id [19] & ((\Mux35~16_combout  & ((\Mux35~18_combout ))) # (!\Mux35~16_combout  & (\Mux35~11_combout )))) # (!\prif.imemload_id [19] & (((\Mux35~16_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\Mux35~11_combout ),
	.datac(\Mux35~18_combout ),
	.datad(\Mux35~16_combout ),
	.cin(gnd),
	.combout(Mux351),
	.cout());
// synopsys translate_off
defparam \Mux35~19 .lut_mask = 16'hF588;
defparam \Mux35~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N26
cycloneive_lcell_comb \Mux37~9 (
// Equation(s):
// Mux37 = (\Mux37~6_combout  & (((\Mux37~8_combout ) # (!\prif.imemload_id [16])))) # (!\Mux37~6_combout  & (\Mux37~1_combout  & (\prif.imemload_id [16])))

	.dataa(\Mux37~6_combout ),
	.datab(\Mux37~1_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux37~8_combout ),
	.cin(gnd),
	.combout(Mux37),
	.cout());
// synopsys translate_off
defparam \Mux37~9 .lut_mask = 16'hEA4A;
defparam \Mux37~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N0
cycloneive_lcell_comb \Mux37~19 (
// Equation(s):
// Mux371 = (\prif.imemload_id [19] & ((\Mux37~16_combout  & ((\Mux37~18_combout ))) # (!\Mux37~16_combout  & (\Mux37~11_combout )))) # (!\prif.imemload_id [19] & (((\Mux37~16_combout ))))

	.dataa(\Mux37~11_combout ),
	.datab(prifimemload_id_19),
	.datac(\Mux37~18_combout ),
	.datad(\Mux37~16_combout ),
	.cin(gnd),
	.combout(Mux371),
	.cout());
// synopsys translate_off
defparam \Mux37~19 .lut_mask = 16'hF388;
defparam \Mux37~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N6
cycloneive_lcell_comb \Mux55~9 (
// Equation(s):
// Mux55 = (\prif.imemload_id [16] & ((\Mux55~6_combout  & ((\Mux55~8_combout ))) # (!\Mux55~6_combout  & (\Mux55~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux55~6_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\Mux55~1_combout ),
	.datac(\Mux55~8_combout ),
	.datad(\Mux55~6_combout ),
	.cin(gnd),
	.combout(Mux55),
	.cout());
// synopsys translate_off
defparam \Mux55~9 .lut_mask = 16'hF588;
defparam \Mux55~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N26
cycloneive_lcell_comb \Mux55~19 (
// Equation(s):
// Mux551 = (\Mux55~16_combout  & (((\Mux55~18_combout )) # (!\prif.imemload_id [19]))) # (!\Mux55~16_combout  & (\prif.imemload_id [19] & (\Mux55~11_combout )))

	.dataa(\Mux55~16_combout ),
	.datab(prifimemload_id_19),
	.datac(\Mux55~11_combout ),
	.datad(\Mux55~18_combout ),
	.cin(gnd),
	.combout(Mux551),
	.cout());
// synopsys translate_off
defparam \Mux55~19 .lut_mask = 16'hEA62;
defparam \Mux55~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N2
cycloneive_lcell_comb \Mux56~9 (
// Equation(s):
// Mux56 = (\prif.imemload_id [16] & ((\Mux56~6_combout  & (\Mux56~8_combout )) # (!\Mux56~6_combout  & ((\Mux56~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux56~6_combout ))))

	.dataa(\Mux56~8_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux56~1_combout ),
	.datad(\Mux56~6_combout ),
	.cin(gnd),
	.combout(Mux56),
	.cout());
// synopsys translate_off
defparam \Mux56~9 .lut_mask = 16'hBBC0;
defparam \Mux56~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N22
cycloneive_lcell_comb \Mux56~19 (
// Equation(s):
// Mux561 = (\prif.imemload_id [18] & ((\Mux56~16_combout  & ((\Mux56~18_combout ))) # (!\Mux56~16_combout  & (\Mux56~11_combout )))) # (!\prif.imemload_id [18] & (((\Mux56~16_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux56~11_combout ),
	.datac(\Mux56~18_combout ),
	.datad(\Mux56~16_combout ),
	.cin(gnd),
	.combout(Mux561),
	.cout());
// synopsys translate_off
defparam \Mux56~19 .lut_mask = 16'hF588;
defparam \Mux56~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N26
cycloneive_lcell_comb \Mux41~9 (
// Equation(s):
// Mux41 = (\prif.imemload_id [16] & ((\Mux41~6_combout  & ((\Mux41~8_combout ))) # (!\Mux41~6_combout  & (\Mux41~1_combout )))) # (!\prif.imemload_id [16] & (((\Mux41~6_combout ))))

	.dataa(\Mux41~1_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux41~8_combout ),
	.datad(\Mux41~6_combout ),
	.cin(gnd),
	.combout(Mux41),
	.cout());
// synopsys translate_off
defparam \Mux41~9 .lut_mask = 16'hF388;
defparam \Mux41~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N14
cycloneive_lcell_comb \Mux41~19 (
// Equation(s):
// Mux411 = (\prif.imemload_id [19] & ((\Mux41~16_combout  & (\Mux41~18_combout )) # (!\Mux41~16_combout  & ((\Mux41~11_combout ))))) # (!\prif.imemload_id [19] & (((\Mux41~16_combout ))))

	.dataa(\Mux41~18_combout ),
	.datab(\Mux41~11_combout ),
	.datac(prifimemload_id_19),
	.datad(\Mux41~16_combout ),
	.cin(gnd),
	.combout(Mux411),
	.cout());
// synopsys translate_off
defparam \Mux41~19 .lut_mask = 16'hAFC0;
defparam \Mux41~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N6
cycloneive_lcell_comb \Mux38~9 (
// Equation(s):
// Mux38 = (\prif.imemload_id [16] & ((\Mux38~6_combout  & (\Mux38~8_combout )) # (!\Mux38~6_combout  & ((\Mux38~1_combout ))))) # (!\prif.imemload_id [16] & (((\Mux38~6_combout ))))

	.dataa(\Mux38~8_combout ),
	.datab(prifimemload_id_16),
	.datac(\Mux38~1_combout ),
	.datad(\Mux38~6_combout ),
	.cin(gnd),
	.combout(Mux38),
	.cout());
// synopsys translate_off
defparam \Mux38~9 .lut_mask = 16'hBBC0;
defparam \Mux38~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N24
cycloneive_lcell_comb \Mux38~19 (
// Equation(s):
// Mux381 = (\Mux38~16_combout  & ((\Mux38~18_combout ) # ((!\prif.imemload_id [18])))) # (!\Mux38~16_combout  & (((\prif.imemload_id [18] & \Mux38~11_combout ))))

	.dataa(\Mux38~18_combout ),
	.datab(\Mux38~16_combout ),
	.datac(prifimemload_id_18),
	.datad(\Mux38~11_combout ),
	.cin(gnd),
	.combout(Mux381),
	.cout());
// synopsys translate_off
defparam \Mux38~19 .lut_mask = 16'hBC8C;
defparam \Mux38~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N16
cycloneive_lcell_comb \Mux29~9 (
// Equation(s):
// Mux29 = (\prif.imemload_id [21] & ((\Mux29~6_combout  & ((\Mux29~8_combout ))) # (!\Mux29~6_combout  & (\Mux29~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux29~6_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\Mux29~1_combout ),
	.datac(\Mux29~8_combout ),
	.datad(\Mux29~6_combout ),
	.cin(gnd),
	.combout(Mux29),
	.cout());
// synopsys translate_off
defparam \Mux29~9 .lut_mask = 16'hF588;
defparam \Mux29~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N4
cycloneive_lcell_comb \Mux29~19 (
// Equation(s):
// Mux291 = (\prif.imemload_id [23] & ((\Mux29~16_combout  & (\Mux29~18_combout )) # (!\Mux29~16_combout  & ((\Mux29~11_combout ))))) # (!\prif.imemload_id [23] & (((\Mux29~16_combout ))))

	.dataa(\Mux29~18_combout ),
	.datab(\Mux29~11_combout ),
	.datac(prifimemload_id_23),
	.datad(\Mux29~16_combout ),
	.cin(gnd),
	.combout(Mux291),
	.cout());
// synopsys translate_off
defparam \Mux29~19 .lut_mask = 16'hAFC0;
defparam \Mux29~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N20
cycloneive_lcell_comb \Mux27~9 (
// Equation(s):
// Mux27 = (\prif.imemload_id [21] & ((\Mux27~6_combout  & ((\Mux27~8_combout ))) # (!\Mux27~6_combout  & (\Mux27~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux27~6_combout ))))

	.dataa(\Mux27~1_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux27~8_combout ),
	.datad(\Mux27~6_combout ),
	.cin(gnd),
	.combout(Mux27),
	.cout());
// synopsys translate_off
defparam \Mux27~9 .lut_mask = 16'hF388;
defparam \Mux27~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N22
cycloneive_lcell_comb \Mux27~19 (
// Equation(s):
// Mux271 = (\prif.imemload_id [23] & ((\Mux27~16_combout  & ((\Mux27~18_combout ))) # (!\Mux27~16_combout  & (\Mux27~11_combout )))) # (!\prif.imemload_id [23] & (((\Mux27~16_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\Mux27~11_combout ),
	.datac(\Mux27~18_combout ),
	.datad(\Mux27~16_combout ),
	.cin(gnd),
	.combout(Mux271),
	.cout());
// synopsys translate_off
defparam \Mux27~19 .lut_mask = 16'hF588;
defparam \Mux27~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N2
cycloneive_lcell_comb \Mux28~9 (
// Equation(s):
// Mux28 = (\prif.imemload_id [21] & ((\Mux28~6_combout  & (\Mux28~8_combout )) # (!\Mux28~6_combout  & ((\Mux28~1_combout ))))) # (!\prif.imemload_id [21] & (((\Mux28~6_combout ))))

	.dataa(\Mux28~8_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux28~6_combout ),
	.datad(\Mux28~1_combout ),
	.cin(gnd),
	.combout(Mux28),
	.cout());
// synopsys translate_off
defparam \Mux28~9 .lut_mask = 16'hBCB0;
defparam \Mux28~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N20
cycloneive_lcell_comb \Mux28~19 (
// Equation(s):
// Mux281 = (\prif.imemload_id [24] & ((\Mux28~16_combout  & ((\Mux28~18_combout ))) # (!\Mux28~16_combout  & (\Mux28~11_combout )))) # (!\prif.imemload_id [24] & (\Mux28~16_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux28~16_combout ),
	.datac(\Mux28~11_combout ),
	.datad(\Mux28~18_combout ),
	.cin(gnd),
	.combout(Mux281),
	.cout());
// synopsys translate_off
defparam \Mux28~19 .lut_mask = 16'hEC64;
defparam \Mux28~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N28
cycloneive_lcell_comb \Mux23~9 (
// Equation(s):
// Mux23 = (\prif.imemload_id [21] & ((\Mux23~6_combout  & (\Mux23~8_combout )) # (!\Mux23~6_combout  & ((\Mux23~1_combout ))))) # (!\prif.imemload_id [21] & (((\Mux23~6_combout ))))

	.dataa(\Mux23~8_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux23~6_combout ),
	.datad(\Mux23~1_combout ),
	.cin(gnd),
	.combout(Mux23),
	.cout());
// synopsys translate_off
defparam \Mux23~9 .lut_mask = 16'hBCB0;
defparam \Mux23~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N6
cycloneive_lcell_comb \Mux23~19 (
// Equation(s):
// Mux231 = (\prif.imemload_id [23] & ((\Mux23~16_combout  & ((\Mux23~18_combout ))) # (!\Mux23~16_combout  & (\Mux23~11_combout )))) # (!\prif.imemload_id [23] & (((\Mux23~16_combout ))))

	.dataa(\Mux23~11_combout ),
	.datab(prifimemload_id_23),
	.datac(\Mux23~18_combout ),
	.datad(\Mux23~16_combout ),
	.cin(gnd),
	.combout(Mux231),
	.cout());
// synopsys translate_off
defparam \Mux23~19 .lut_mask = 16'hF388;
defparam \Mux23~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N18
cycloneive_lcell_comb \Mux24~9 (
// Equation(s):
// Mux24 = (\Mux24~6_combout  & ((\Mux24~8_combout ) # ((!\prif.imemload_id [21])))) # (!\Mux24~6_combout  & (((\prif.imemload_id [21] & \Mux24~1_combout ))))

	.dataa(\Mux24~8_combout ),
	.datab(\Mux24~6_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux24~1_combout ),
	.cin(gnd),
	.combout(Mux24),
	.cout());
// synopsys translate_off
defparam \Mux24~9 .lut_mask = 16'hBC8C;
defparam \Mux24~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N4
cycloneive_lcell_comb \Mux24~19 (
// Equation(s):
// Mux241 = (\prif.imemload_id [24] & ((\Mux24~16_combout  & (\Mux24~18_combout )) # (!\Mux24~16_combout  & ((\Mux24~11_combout ))))) # (!\prif.imemload_id [24] & (((\Mux24~16_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\Mux24~18_combout ),
	.datac(\Mux24~11_combout ),
	.datad(\Mux24~16_combout ),
	.cin(gnd),
	.combout(Mux241),
	.cout());
// synopsys translate_off
defparam \Mux24~19 .lut_mask = 16'hDDA0;
defparam \Mux24~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N26
cycloneive_lcell_comb \Mux25~9 (
// Equation(s):
// Mux25 = (\Mux25~6_combout  & ((\Mux25~8_combout ) # ((!\prif.imemload_id [21])))) # (!\Mux25~6_combout  & (((\prif.imemload_id [21] & \Mux25~1_combout ))))

	.dataa(\Mux25~8_combout ),
	.datab(\Mux25~6_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux25~1_combout ),
	.cin(gnd),
	.combout(Mux25),
	.cout());
// synopsys translate_off
defparam \Mux25~9 .lut_mask = 16'hBC8C;
defparam \Mux25~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N20
cycloneive_lcell_comb \Mux25~19 (
// Equation(s):
// Mux251 = (\Mux25~16_combout  & ((\Mux25~18_combout ) # ((!\prif.imemload_id [23])))) # (!\Mux25~16_combout  & (((\prif.imemload_id [23] & \Mux25~11_combout ))))

	.dataa(\Mux25~18_combout ),
	.datab(\Mux25~16_combout ),
	.datac(prifimemload_id_23),
	.datad(\Mux25~11_combout ),
	.cin(gnd),
	.combout(Mux251),
	.cout());
// synopsys translate_off
defparam \Mux25~19 .lut_mask = 16'hBC8C;
defparam \Mux25~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N28
cycloneive_lcell_comb \Mux26~9 (
// Equation(s):
// Mux26 = (\Mux26~6_combout  & (((\Mux26~8_combout ) # (!\prif.imemload_id [21])))) # (!\Mux26~6_combout  & (\Mux26~1_combout  & ((\prif.imemload_id [21]))))

	.dataa(\Mux26~1_combout ),
	.datab(\Mux26~8_combout ),
	.datac(\Mux26~6_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(Mux26),
	.cout());
// synopsys translate_off
defparam \Mux26~9 .lut_mask = 16'hCAF0;
defparam \Mux26~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N14
cycloneive_lcell_comb \Mux26~19 (
// Equation(s):
// Mux261 = (\Mux26~16_combout  & ((\Mux26~18_combout ) # ((!\prif.imemload_id [24])))) # (!\Mux26~16_combout  & (((\prif.imemload_id [24] & \Mux26~11_combout ))))

	.dataa(\Mux26~16_combout ),
	.datab(\Mux26~18_combout ),
	.datac(prifimemload_id_24),
	.datad(\Mux26~11_combout ),
	.cin(gnd),
	.combout(Mux261),
	.cout());
// synopsys translate_off
defparam \Mux26~19 .lut_mask = 16'hDA8A;
defparam \Mux26~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N16
cycloneive_lcell_comb \Mux15~9 (
// Equation(s):
// Mux15 = (\prif.imemload_id [21] & ((\Mux15~6_combout  & (\Mux15~8_combout )) # (!\Mux15~6_combout  & ((\Mux15~1_combout ))))) # (!\prif.imemload_id [21] & (((\Mux15~6_combout ))))

	.dataa(\Mux15~8_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux15~1_combout ),
	.datad(\Mux15~6_combout ),
	.cin(gnd),
	.combout(Mux15),
	.cout());
// synopsys translate_off
defparam \Mux15~9 .lut_mask = 16'hBBC0;
defparam \Mux15~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N28
cycloneive_lcell_comb \Mux15~19 (
// Equation(s):
// Mux1510 = (\prif.imemload_id [23] & ((\Mux15~16_combout  & (\Mux15~18_combout )) # (!\Mux15~16_combout  & ((\Mux15~11_combout ))))) # (!\prif.imemload_id [23] & (((\Mux15~16_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\Mux15~18_combout ),
	.datac(\Mux15~16_combout ),
	.datad(\Mux15~11_combout ),
	.cin(gnd),
	.combout(Mux1510),
	.cout());
// synopsys translate_off
defparam \Mux15~19 .lut_mask = 16'hDAD0;
defparam \Mux15~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y24_N2
cycloneive_lcell_comb \Mux16~9 (
// Equation(s):
// Mux16 = (\prif.imemload_id [21] & ((\Mux16~6_combout  & ((\Mux16~8_combout ))) # (!\Mux16~6_combout  & (\Mux16~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux16~6_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\Mux16~1_combout ),
	.datac(\Mux16~8_combout ),
	.datad(\Mux16~6_combout ),
	.cin(gnd),
	.combout(Mux16),
	.cout());
// synopsys translate_off
defparam \Mux16~9 .lut_mask = 16'hF588;
defparam \Mux16~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N22
cycloneive_lcell_comb \Mux16~19 (
// Equation(s):
// Mux165 = (\prif.imemload_id [24] & ((\Mux16~16_combout  & (\Mux16~18_combout )) # (!\Mux16~16_combout  & ((\Mux16~11_combout ))))) # (!\prif.imemload_id [24] & (((\Mux16~16_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\Mux16~18_combout ),
	.datac(\Mux16~11_combout ),
	.datad(\Mux16~16_combout ),
	.cin(gnd),
	.combout(Mux165),
	.cout());
// synopsys translate_off
defparam \Mux16~19 .lut_mask = 16'hDDA0;
defparam \Mux16~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N18
cycloneive_lcell_comb \Mux17~9 (
// Equation(s):
// Mux17 = (\prif.imemload_id [21] & ((\Mux17~6_combout  & ((\Mux17~8_combout ))) # (!\Mux17~6_combout  & (\Mux17~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux17~6_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\Mux17~1_combout ),
	.datac(\Mux17~8_combout ),
	.datad(\Mux17~6_combout ),
	.cin(gnd),
	.combout(Mux17),
	.cout());
// synopsys translate_off
defparam \Mux17~9 .lut_mask = 16'hF588;
defparam \Mux17~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N30
cycloneive_lcell_comb \Mux17~19 (
// Equation(s):
// Mux171 = (\prif.imemload_id [23] & ((\Mux17~16_combout  & (\Mux17~18_combout )) # (!\Mux17~16_combout  & ((\Mux17~11_combout ))))) # (!\prif.imemload_id [23] & (\Mux17~16_combout ))

	.dataa(prifimemload_id_23),
	.datab(\Mux17~16_combout ),
	.datac(\Mux17~18_combout ),
	.datad(\Mux17~11_combout ),
	.cin(gnd),
	.combout(Mux171),
	.cout());
// synopsys translate_off
defparam \Mux17~19 .lut_mask = 16'hE6C4;
defparam \Mux17~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N12
cycloneive_lcell_comb \Mux18~9 (
// Equation(s):
// Mux18 = (\prif.imemload_id [21] & ((\Mux18~6_combout  & ((\Mux18~8_combout ))) # (!\Mux18~6_combout  & (\Mux18~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux18~6_combout ))))

	.dataa(\Mux18~1_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux18~8_combout ),
	.datad(\Mux18~6_combout ),
	.cin(gnd),
	.combout(Mux18),
	.cout());
// synopsys translate_off
defparam \Mux18~9 .lut_mask = 16'hF388;
defparam \Mux18~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N22
cycloneive_lcell_comb \Mux18~19 (
// Equation(s):
// Mux181 = (\prif.imemload_id [24] & ((\Mux18~16_combout  & (\Mux18~18_combout )) # (!\Mux18~16_combout  & ((\Mux18~11_combout ))))) # (!\prif.imemload_id [24] & (((\Mux18~16_combout ))))

	.dataa(\Mux18~18_combout ),
	.datab(\Mux18~11_combout ),
	.datac(prifimemload_id_24),
	.datad(\Mux18~16_combout ),
	.cin(gnd),
	.combout(Mux181),
	.cout());
// synopsys translate_off
defparam \Mux18~19 .lut_mask = 16'hAFC0;
defparam \Mux18~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N8
cycloneive_lcell_comb \Mux20~9 (
// Equation(s):
// Mux20 = (\prif.imemload_id [21] & ((\Mux20~6_combout  & ((\Mux20~8_combout ))) # (!\Mux20~6_combout  & (\Mux20~1_combout )))) # (!\prif.imemload_id [21] & (\Mux20~6_combout ))

	.dataa(prifimemload_id_21),
	.datab(\Mux20~6_combout ),
	.datac(\Mux20~1_combout ),
	.datad(\Mux20~8_combout ),
	.cin(gnd),
	.combout(Mux20),
	.cout());
// synopsys translate_off
defparam \Mux20~9 .lut_mask = 16'hEC64;
defparam \Mux20~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N2
cycloneive_lcell_comb \Mux20~19 (
// Equation(s):
// Mux201 = (\prif.imemload_id [24] & ((\Mux20~16_combout  & ((\Mux20~18_combout ))) # (!\Mux20~16_combout  & (\Mux20~11_combout )))) # (!\prif.imemload_id [24] & (\Mux20~16_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux20~16_combout ),
	.datac(\Mux20~11_combout ),
	.datad(\Mux20~18_combout ),
	.cin(gnd),
	.combout(Mux201),
	.cout());
// synopsys translate_off
defparam \Mux20~19 .lut_mask = 16'hEC64;
defparam \Mux20~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N28
cycloneive_lcell_comb \Mux19~9 (
// Equation(s):
// Mux19 = (\prif.imemload_id [21] & ((\Mux19~6_combout  & (\Mux19~8_combout )) # (!\Mux19~6_combout  & ((\Mux19~1_combout ))))) # (!\prif.imemload_id [21] & (((\Mux19~6_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\Mux19~8_combout ),
	.datac(\Mux19~1_combout ),
	.datad(\Mux19~6_combout ),
	.cin(gnd),
	.combout(Mux19),
	.cout());
// synopsys translate_off
defparam \Mux19~9 .lut_mask = 16'hDDA0;
defparam \Mux19~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N0
cycloneive_lcell_comb \Mux19~19 (
// Equation(s):
// Mux191 = (\prif.imemload_id [23] & ((\Mux19~16_combout  & ((\Mux19~18_combout ))) # (!\Mux19~16_combout  & (\Mux19~11_combout )))) # (!\prif.imemload_id [23] & (((\Mux19~16_combout ))))

	.dataa(\Mux19~11_combout ),
	.datab(\Mux19~18_combout ),
	.datac(prifimemload_id_23),
	.datad(\Mux19~16_combout ),
	.cin(gnd),
	.combout(Mux191),
	.cout());
// synopsys translate_off
defparam \Mux19~19 .lut_mask = 16'hCFA0;
defparam \Mux19~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N2
cycloneive_lcell_comb \Mux21~9 (
// Equation(s):
// Mux21 = (\Mux21~6_combout  & ((\Mux21~8_combout ) # ((!\prif.imemload_id [21])))) # (!\Mux21~6_combout  & (((\Mux21~1_combout  & \prif.imemload_id [21]))))

	.dataa(\Mux21~8_combout ),
	.datab(\Mux21~6_combout ),
	.datac(\Mux21~1_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(Mux21),
	.cout());
// synopsys translate_off
defparam \Mux21~9 .lut_mask = 16'hB8CC;
defparam \Mux21~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N26
cycloneive_lcell_comb \Mux21~19 (
// Equation(s):
// Mux211 = (\prif.imemload_id [23] & ((\Mux21~16_combout  & ((\Mux21~18_combout ))) # (!\Mux21~16_combout  & (\Mux21~11_combout )))) # (!\prif.imemload_id [23] & (((\Mux21~16_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\Mux21~11_combout ),
	.datac(\Mux21~18_combout ),
	.datad(\Mux21~16_combout ),
	.cin(gnd),
	.combout(Mux211),
	.cout());
// synopsys translate_off
defparam \Mux21~19 .lut_mask = 16'hF588;
defparam \Mux21~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N10
cycloneive_lcell_comb \Mux22~9 (
// Equation(s):
// Mux22 = (\Mux22~6_combout  & (((\Mux22~8_combout ) # (!\prif.imemload_id [21])))) # (!\Mux22~6_combout  & (\Mux22~1_combout  & ((\prif.imemload_id [21]))))

	.dataa(\Mux22~1_combout ),
	.datab(\Mux22~8_combout ),
	.datac(\Mux22~6_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(Mux22),
	.cout());
// synopsys translate_off
defparam \Mux22~9 .lut_mask = 16'hCAF0;
defparam \Mux22~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N16
cycloneive_lcell_comb \Mux22~19 (
// Equation(s):
// Mux221 = (\prif.imemload_id [24] & ((\Mux22~16_combout  & (\Mux22~18_combout )) # (!\Mux22~16_combout  & ((\Mux22~11_combout ))))) # (!\prif.imemload_id [24] & (((\Mux22~16_combout ))))

	.dataa(\Mux22~18_combout ),
	.datab(prifimemload_id_24),
	.datac(\Mux22~11_combout ),
	.datad(\Mux22~16_combout ),
	.cin(gnd),
	.combout(Mux221),
	.cout());
// synopsys translate_off
defparam \Mux22~19 .lut_mask = 16'hBBC0;
defparam \Mux22~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N0
cycloneive_lcell_comb \Mux13~9 (
// Equation(s):
// Mux13 = (\Mux13~6_combout  & ((\Mux13~8_combout ) # ((!\prif.imemload_id [21])))) # (!\Mux13~6_combout  & (((\Mux13~1_combout  & \prif.imemload_id [21]))))

	.dataa(\Mux13~8_combout ),
	.datab(\Mux13~1_combout ),
	.datac(\Mux13~6_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(Mux13),
	.cout());
// synopsys translate_off
defparam \Mux13~9 .lut_mask = 16'hACF0;
defparam \Mux13~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N26
cycloneive_lcell_comb \Mux13~19 (
// Equation(s):
// Mux131 = (\prif.imemload_id [23] & ((\Mux13~16_combout  & ((\Mux13~18_combout ))) # (!\Mux13~16_combout  & (\Mux13~11_combout )))) # (!\prif.imemload_id [23] & (((\Mux13~16_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\Mux13~11_combout ),
	.datac(\Mux13~18_combout ),
	.datad(\Mux13~16_combout ),
	.cin(gnd),
	.combout(Mux131),
	.cout());
// synopsys translate_off
defparam \Mux13~19 .lut_mask = 16'hF588;
defparam \Mux13~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N4
cycloneive_lcell_comb \Mux14~9 (
// Equation(s):
// Mux14 = (\Mux14~6_combout  & (((\Mux14~8_combout ) # (!\prif.imemload_id [21])))) # (!\Mux14~6_combout  & (\Mux14~1_combout  & ((\prif.imemload_id [21]))))

	.dataa(\Mux14~1_combout ),
	.datab(\Mux14~6_combout ),
	.datac(\Mux14~8_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(Mux14),
	.cout());
// synopsys translate_off
defparam \Mux14~9 .lut_mask = 16'hE2CC;
defparam \Mux14~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N30
cycloneive_lcell_comb \Mux14~19 (
// Equation(s):
// Mux1410 = (\Mux14~16_combout  & ((\Mux14~18_combout ) # ((!\prif.imemload_id [24])))) # (!\Mux14~16_combout  & (((\prif.imemload_id [24] & \Mux14~11_combout ))))

	.dataa(\Mux14~18_combout ),
	.datab(\Mux14~16_combout ),
	.datac(prifimemload_id_24),
	.datad(\Mux14~11_combout ),
	.cin(gnd),
	.combout(Mux1410),
	.cout());
// synopsys translate_off
defparam \Mux14~19 .lut_mask = 16'hBC8C;
defparam \Mux14~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N0
cycloneive_lcell_comb \Mux11~9 (
// Equation(s):
// Mux11 = (\prif.imemload_id [21] & ((\Mux11~6_combout  & ((\Mux11~8_combout ))) # (!\Mux11~6_combout  & (\Mux11~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux11~6_combout ))))

	.dataa(\Mux11~1_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux11~8_combout ),
	.datad(\Mux11~6_combout ),
	.cin(gnd),
	.combout(Mux11),
	.cout());
// synopsys translate_off
defparam \Mux11~9 .lut_mask = 16'hF388;
defparam \Mux11~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N22
cycloneive_lcell_comb \Mux11~19 (
// Equation(s):
// Mux111 = (\prif.imemload_id [23] & ((\Mux11~16_combout  & (\Mux11~18_combout )) # (!\Mux11~16_combout  & ((\Mux11~11_combout ))))) # (!\prif.imemload_id [23] & (((\Mux11~16_combout ))))

	.dataa(\Mux11~18_combout ),
	.datab(\Mux11~11_combout ),
	.datac(prifimemload_id_23),
	.datad(\Mux11~16_combout ),
	.cin(gnd),
	.combout(Mux111),
	.cout());
// synopsys translate_off
defparam \Mux11~19 .lut_mask = 16'hAFC0;
defparam \Mux11~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N2
cycloneive_lcell_comb \Mux12~9 (
// Equation(s):
// Mux12 = (\prif.imemload_id [21] & ((\Mux12~6_combout  & ((\Mux12~8_combout ))) # (!\Mux12~6_combout  & (\Mux12~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux12~6_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\Mux12~1_combout ),
	.datac(\Mux12~6_combout ),
	.datad(\Mux12~8_combout ),
	.cin(gnd),
	.combout(Mux12),
	.cout());
// synopsys translate_off
defparam \Mux12~9 .lut_mask = 16'hF858;
defparam \Mux12~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N8
cycloneive_lcell_comb \Mux12~19 (
// Equation(s):
// Mux121 = (\prif.imemload_id [24] & ((\Mux12~16_combout  & ((\Mux12~18_combout ))) # (!\Mux12~16_combout  & (\Mux12~11_combout )))) # (!\prif.imemload_id [24] & (((\Mux12~16_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\Mux12~11_combout ),
	.datac(\Mux12~18_combout ),
	.datad(\Mux12~16_combout ),
	.cin(gnd),
	.combout(Mux121),
	.cout());
// synopsys translate_off
defparam \Mux12~19 .lut_mask = 16'hF588;
defparam \Mux12~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N30
cycloneive_lcell_comb \Mux9~9 (
// Equation(s):
// Mux9 = (\Mux9~6_combout  & (((\Mux9~8_combout ) # (!\prif.imemload_id [21])))) # (!\Mux9~6_combout  & (\Mux9~1_combout  & ((\prif.imemload_id [21]))))

	.dataa(\Mux9~1_combout ),
	.datab(\Mux9~8_combout ),
	.datac(\Mux9~6_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(Mux9),
	.cout());
// synopsys translate_off
defparam \Mux9~9 .lut_mask = 16'hCAF0;
defparam \Mux9~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N14
cycloneive_lcell_comb \Mux9~19 (
// Equation(s):
// Mux91 = (\prif.imemload_id [23] & ((\Mux9~16_combout  & (\Mux9~18_combout )) # (!\Mux9~16_combout  & ((\Mux9~11_combout ))))) # (!\prif.imemload_id [23] & (((\Mux9~16_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\Mux9~18_combout ),
	.datac(\Mux9~11_combout ),
	.datad(\Mux9~16_combout ),
	.cin(gnd),
	.combout(Mux91),
	.cout());
// synopsys translate_off
defparam \Mux9~19 .lut_mask = 16'hDDA0;
defparam \Mux9~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N24
cycloneive_lcell_comb \Mux10~9 (
// Equation(s):
// Mux10 = (\Mux10~6_combout  & ((\Mux10~8_combout ) # ((!\prif.imemload_id [21])))) # (!\Mux10~6_combout  & (((\prif.imemload_id [21] & \Mux10~1_combout ))))

	.dataa(\Mux10~6_combout ),
	.datab(\Mux10~8_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux10~1_combout ),
	.cin(gnd),
	.combout(Mux10),
	.cout());
// synopsys translate_off
defparam \Mux10~9 .lut_mask = 16'hDA8A;
defparam \Mux10~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N4
cycloneive_lcell_comb \Mux10~19 (
// Equation(s):
// Mux101 = (\prif.imemload_id [24] & ((\Mux10~16_combout  & ((\Mux10~18_combout ))) # (!\Mux10~16_combout  & (\Mux10~11_combout )))) # (!\prif.imemload_id [24] & (((\Mux10~16_combout ))))

	.dataa(\Mux10~11_combout ),
	.datab(\Mux10~18_combout ),
	.datac(prifimemload_id_24),
	.datad(\Mux10~16_combout ),
	.cin(gnd),
	.combout(Mux101),
	.cout());
// synopsys translate_off
defparam \Mux10~19 .lut_mask = 16'hCFA0;
defparam \Mux10~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N30
cycloneive_lcell_comb \Mux7~9 (
// Equation(s):
// Mux7 = (\prif.imemload_id [21] & ((\Mux7~6_combout  & (\Mux7~8_combout )) # (!\Mux7~6_combout  & ((\Mux7~1_combout ))))) # (!\prif.imemload_id [21] & (((\Mux7~6_combout ))))

	.dataa(\Mux7~8_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux7~1_combout ),
	.datad(\Mux7~6_combout ),
	.cin(gnd),
	.combout(Mux7),
	.cout());
// synopsys translate_off
defparam \Mux7~9 .lut_mask = 16'hBBC0;
defparam \Mux7~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N24
cycloneive_lcell_comb \Mux7~19 (
// Equation(s):
// Mux71 = (\prif.imemload_id [23] & ((\Mux7~16_combout  & (\Mux7~18_combout )) # (!\Mux7~16_combout  & ((\Mux7~11_combout ))))) # (!\prif.imemload_id [23] & (((\Mux7~16_combout ))))

	.dataa(\Mux7~18_combout ),
	.datab(prifimemload_id_23),
	.datac(\Mux7~11_combout ),
	.datad(\Mux7~16_combout ),
	.cin(gnd),
	.combout(Mux71),
	.cout());
// synopsys translate_off
defparam \Mux7~19 .lut_mask = 16'hBBC0;
defparam \Mux7~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N10
cycloneive_lcell_comb \Mux8~9 (
// Equation(s):
// Mux8 = (\prif.imemload_id [21] & ((\Mux8~6_combout  & ((\Mux8~8_combout ))) # (!\Mux8~6_combout  & (\Mux8~1_combout )))) # (!\prif.imemload_id [21] & (\Mux8~6_combout ))

	.dataa(prifimemload_id_21),
	.datab(\Mux8~6_combout ),
	.datac(\Mux8~1_combout ),
	.datad(\Mux8~8_combout ),
	.cin(gnd),
	.combout(Mux8),
	.cout());
// synopsys translate_off
defparam \Mux8~9 .lut_mask = 16'hEC64;
defparam \Mux8~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N18
cycloneive_lcell_comb \Mux8~19 (
// Equation(s):
// Mux81 = (\prif.imemload_id [24] & ((\Mux8~16_combout  & ((\Mux8~18_combout ))) # (!\Mux8~16_combout  & (\Mux8~11_combout )))) # (!\prif.imemload_id [24] & (\Mux8~16_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux8~16_combout ),
	.datac(\Mux8~11_combout ),
	.datad(\Mux8~18_combout ),
	.cin(gnd),
	.combout(Mux81),
	.cout());
// synopsys translate_off
defparam \Mux8~19 .lut_mask = 16'hEC64;
defparam \Mux8~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N8
cycloneive_lcell_comb \Mux0~9 (
// Equation(s):
// Mux0 = (\prif.imemload_id [21] & ((\Mux0~6_combout  & ((\Mux0~8_combout ))) # (!\Mux0~6_combout  & (\Mux0~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux0~6_combout ))))

	.dataa(\Mux0~1_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux0~8_combout ),
	.datad(\Mux0~6_combout ),
	.cin(gnd),
	.combout(Mux0),
	.cout());
// synopsys translate_off
defparam \Mux0~9 .lut_mask = 16'hF388;
defparam \Mux0~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N24
cycloneive_lcell_comb \Mux0~19 (
// Equation(s):
// Mux01 = (\prif.imemload_id [24] & ((\Mux0~16_combout  & (\Mux0~18_combout )) # (!\Mux0~16_combout  & ((\Mux0~11_combout ))))) # (!\prif.imemload_id [24] & (((\Mux0~16_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\Mux0~18_combout ),
	.datac(\Mux0~11_combout ),
	.datad(\Mux0~16_combout ),
	.cin(gnd),
	.combout(Mux01),
	.cout());
// synopsys translate_off
defparam \Mux0~19 .lut_mask = 16'hDDA0;
defparam \Mux0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N0
cycloneive_lcell_comb \Mux1~9 (
// Equation(s):
// Mux1 = (\prif.imemload_id [21] & ((\Mux1~6_combout  & ((\Mux1~8_combout ))) # (!\Mux1~6_combout  & (\Mux1~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux1~6_combout ))))

	.dataa(\Mux1~1_combout ),
	.datab(\Mux1~8_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux1~6_combout ),
	.cin(gnd),
	.combout(Mux1),
	.cout());
// synopsys translate_off
defparam \Mux1~9 .lut_mask = 16'hCFA0;
defparam \Mux1~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N22
cycloneive_lcell_comb \Mux1~19 (
// Equation(s):
// Mux110 = (\prif.imemload_id [23] & ((\Mux1~16_combout  & (\Mux1~18_combout )) # (!\Mux1~16_combout  & ((\Mux1~11_combout ))))) # (!\prif.imemload_id [23] & (((\Mux1~16_combout ))))

	.dataa(\Mux1~18_combout ),
	.datab(prifimemload_id_23),
	.datac(\Mux1~11_combout ),
	.datad(\Mux1~16_combout ),
	.cin(gnd),
	.combout(Mux110),
	.cout());
// synopsys translate_off
defparam \Mux1~19 .lut_mask = 16'hBBC0;
defparam \Mux1~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N28
cycloneive_lcell_comb \Mux2~9 (
// Equation(s):
// Mux2 = (\Mux2~6_combout  & (((\Mux2~8_combout ) # (!\prif.imemload_id [21])))) # (!\Mux2~6_combout  & (\Mux2~1_combout  & (\prif.imemload_id [21])))

	.dataa(\Mux2~6_combout ),
	.datab(\Mux2~1_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux2~8_combout ),
	.cin(gnd),
	.combout(Mux2),
	.cout());
// synopsys translate_off
defparam \Mux2~9 .lut_mask = 16'hEA4A;
defparam \Mux2~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N8
cycloneive_lcell_comb \Mux2~19 (
// Equation(s):
// Mux210 = (\Mux2~16_combout  & ((\Mux2~18_combout ) # ((!\prif.imemload_id [24])))) # (!\Mux2~16_combout  & (((\prif.imemload_id [24] & \Mux2~11_combout ))))

	.dataa(\Mux2~16_combout ),
	.datab(\Mux2~18_combout ),
	.datac(prifimemload_id_24),
	.datad(\Mux2~11_combout ),
	.cin(gnd),
	.combout(Mux210),
	.cout());
// synopsys translate_off
defparam \Mux2~19 .lut_mask = 16'hDA8A;
defparam \Mux2~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N12
cycloneive_lcell_comb \Mux5~9 (
// Equation(s):
// Mux5 = (\prif.imemload_id [21] & ((\Mux5~6_combout  & (\Mux5~8_combout )) # (!\Mux5~6_combout  & ((\Mux5~1_combout ))))) # (!\prif.imemload_id [21] & (((\Mux5~6_combout ))))

	.dataa(\Mux5~8_combout ),
	.datab(\Mux5~1_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux5~6_combout ),
	.cin(gnd),
	.combout(Mux5),
	.cout());
// synopsys translate_off
defparam \Mux5~9 .lut_mask = 16'hAFC0;
defparam \Mux5~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N28
cycloneive_lcell_comb \Mux5~19 (
// Equation(s):
// Mux510 = (\prif.imemload_id [23] & ((\Mux5~16_combout  & (\Mux5~18_combout )) # (!\Mux5~16_combout  & ((\Mux5~11_combout ))))) # (!\prif.imemload_id [23] & (((\Mux5~16_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\Mux5~18_combout ),
	.datac(\Mux5~11_combout ),
	.datad(\Mux5~16_combout ),
	.cin(gnd),
	.combout(Mux510),
	.cout());
// synopsys translate_off
defparam \Mux5~19 .lut_mask = 16'hDDA0;
defparam \Mux5~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N18
cycloneive_lcell_comb \Mux6~9 (
// Equation(s):
// Mux6 = (\prif.imemload_id [21] & ((\Mux6~6_combout  & ((\Mux6~8_combout ))) # (!\Mux6~6_combout  & (\Mux6~1_combout )))) # (!\prif.imemload_id [21] & (((\Mux6~6_combout ))))

	.dataa(\Mux6~1_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux6~8_combout ),
	.datad(\Mux6~6_combout ),
	.cin(gnd),
	.combout(Mux6),
	.cout());
// synopsys translate_off
defparam \Mux6~9 .lut_mask = 16'hF388;
defparam \Mux6~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N24
cycloneive_lcell_comb \Mux6~19 (
// Equation(s):
// Mux64 = (\prif.imemload_id [24] & ((\Mux6~16_combout  & ((\Mux6~18_combout ))) # (!\Mux6~16_combout  & (\Mux6~11_combout )))) # (!\prif.imemload_id [24] & (((\Mux6~16_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\Mux6~11_combout ),
	.datac(\Mux6~16_combout ),
	.datad(\Mux6~18_combout ),
	.cin(gnd),
	.combout(Mux64),
	.cout());
// synopsys translate_off
defparam \Mux6~19 .lut_mask = 16'hF858;
defparam \Mux6~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N6
cycloneive_lcell_comb \Mux3~9 (
// Equation(s):
// Mux3 = (\prif.imemload_id [21] & ((\Mux3~6_combout  & (\Mux3~8_combout )) # (!\Mux3~6_combout  & ((\Mux3~1_combout ))))) # (!\prif.imemload_id [21] & (((\Mux3~6_combout ))))

	.dataa(\Mux3~8_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux3~1_combout ),
	.datad(\Mux3~6_combout ),
	.cin(gnd),
	.combout(Mux3),
	.cout());
// synopsys translate_off
defparam \Mux3~9 .lut_mask = 16'hBBC0;
defparam \Mux3~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N30
cycloneive_lcell_comb \Mux3~19 (
// Equation(s):
// Mux310 = (\prif.imemload_id [23] & ((\Mux3~16_combout  & ((\Mux3~18_combout ))) # (!\Mux3~16_combout  & (\Mux3~11_combout )))) # (!\prif.imemload_id [23] & (((\Mux3~16_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\Mux3~11_combout ),
	.datac(\Mux3~16_combout ),
	.datad(\Mux3~18_combout ),
	.cin(gnd),
	.combout(Mux310),
	.cout());
// synopsys translate_off
defparam \Mux3~19 .lut_mask = 16'hF858;
defparam \Mux3~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N8
cycloneive_lcell_comb \Mux4~9 (
// Equation(s):
// Mux4 = (\Mux4~6_combout  & (((\Mux4~8_combout ) # (!\prif.imemload_id [21])))) # (!\Mux4~6_combout  & (\Mux4~1_combout  & (\prif.imemload_id [21])))

	.dataa(\Mux4~1_combout ),
	.datab(\Mux4~6_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux4~8_combout ),
	.cin(gnd),
	.combout(Mux4),
	.cout());
// synopsys translate_off
defparam \Mux4~9 .lut_mask = 16'hEC2C;
defparam \Mux4~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N12
cycloneive_lcell_comb \Mux4~19 (
// Equation(s):
// Mux410 = (\Mux4~16_combout  & (((\Mux4~18_combout ) # (!\prif.imemload_id [24])))) # (!\Mux4~16_combout  & (\Mux4~11_combout  & ((\prif.imemload_id [24]))))

	.dataa(\Mux4~11_combout ),
	.datab(\Mux4~16_combout ),
	.datac(\Mux4~18_combout ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(Mux410),
	.cout());
// synopsys translate_off
defparam \Mux4~19 .lut_mask = 16'hE2CC;
defparam \Mux4~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N6
cycloneive_lcell_comb \reg_file_nxt[31][1]~64 (
// Equation(s):
// \reg_file_nxt[31][1]~64_combout  = (\Mux163~1_combout  & ((\prif.regwrite_wb [0]) # ((\prif.regwrite_wb [2]) # (!Equal8))))

	.dataa(Mux163),
	.datab(prifregwrite_wb_0),
	.datac(Equal8),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\reg_file_nxt[31][1]~64_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][1]~64 .lut_mask = 16'hAA8A;
defparam \reg_file_nxt[31][1]~64 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N12
cycloneive_lcell_comb \Decoder0~14 (
// Equation(s):
// \Decoder0~14_combout  = (\prif.Regwen_wb~q  & (\prif.regwrite_wb [0] & \prif.regwrite_wb [2]))

	.dataa(prifRegwen_wb),
	.datab(gnd),
	.datac(prifregwrite_wb_0),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\Decoder0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~14 .lut_mask = 16'hA000;
defparam \Decoder0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N26
cycloneive_lcell_comb \Decoder0~15 (
// Equation(s):
// \Decoder0~15_combout  = (!\prif.regwrite_wb [1] & (\prif.regwrite_wb [4] & (\Decoder0~14_combout  & !\prif.regwrite_wb [3])))

	.dataa(prifregwrite_wb_1),
	.datab(prifregwrite_wb_4),
	.datac(\Decoder0~14_combout ),
	.datad(prifregwrite_wb_3),
	.cin(gnd),
	.combout(\Decoder0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~15 .lut_mask = 16'h0040;
defparam \Decoder0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N17
dffeas \reg_file[21][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][1] .is_wysiwyg = "true";
defparam \reg_file[21][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N18
cycloneive_lcell_comb \Decoder0~19 (
// Equation(s):
// \Decoder0~19_combout  = (\prif.regwrite_wb [3] & (\Decoder0~14_combout  & (\prif.regwrite_wb [4] & !\prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~14_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~19_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~19 .lut_mask = 16'h0080;
defparam \Decoder0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N25
dffeas \reg_file[29][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][1] .is_wysiwyg = "true";
defparam \reg_file[29][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N30
cycloneive_lcell_comb \Decoder0~16 (
// Equation(s):
// \Decoder0~16_combout  = (\prif.regwrite_wb [0] & (\prif.Regwen_wb~q  & !\prif.regwrite_wb [2]))

	.dataa(gnd),
	.datab(prifregwrite_wb_0),
	.datac(prifRegwen_wb),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\Decoder0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~16 .lut_mask = 16'h00C0;
defparam \Decoder0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N4
cycloneive_lcell_comb \Decoder0~18 (
// Equation(s):
// \Decoder0~18_combout  = (!\prif.regwrite_wb [1] & (\Decoder0~16_combout  & (\prif.regwrite_wb [4] & !\prif.regwrite_wb [3])))

	.dataa(prifregwrite_wb_1),
	.datab(\Decoder0~16_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_3),
	.cin(gnd),
	.combout(\Decoder0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~18 .lut_mask = 16'h0040;
defparam \Decoder0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N13
dffeas \reg_file[17][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][1] .is_wysiwyg = "true";
defparam \reg_file[17][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N2
cycloneive_lcell_comb \Decoder0~17 (
// Equation(s):
// \Decoder0~17_combout  = (!\prif.regwrite_wb [1] & (\Decoder0~16_combout  & (\prif.regwrite_wb [4] & \prif.regwrite_wb [3])))

	.dataa(prifregwrite_wb_1),
	.datab(\Decoder0~16_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_3),
	.cin(gnd),
	.combout(\Decoder0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~17 .lut_mask = 16'h4000;
defparam \Decoder0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N13
dffeas \reg_file[25][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][1] .is_wysiwyg = "true";
defparam \reg_file[25][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N12
cycloneive_lcell_comb \Mux62~0 (
// Equation(s):
// \Mux62~0_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[25][1]~q ))) # (!\prif.imemload_id [19] & (\reg_file[17][1]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][1]~q ),
	.datad(\reg_file[25][1]~q ),
	.cin(gnd),
	.combout(\Mux62~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~0 .lut_mask = 16'hDC98;
defparam \Mux62~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N24
cycloneive_lcell_comb \Mux62~1 (
// Equation(s):
// \Mux62~1_combout  = (\prif.imemload_id [18] & ((\Mux62~0_combout  & ((\reg_file[29][1]~q ))) # (!\Mux62~0_combout  & (\reg_file[21][1]~q )))) # (!\prif.imemload_id [18] & (((\Mux62~0_combout ))))

	.dataa(\reg_file[21][1]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[29][1]~q ),
	.datad(\Mux62~0_combout ),
	.cin(gnd),
	.combout(\Mux62~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~1 .lut_mask = 16'hF388;
defparam \Mux62~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N24
cycloneive_lcell_comb \reg_file[30][1]~feeder (
// Equation(s):
// \reg_file[30][1]~feeder_combout  = \reg_file_nxt[31][1]~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][1]~64_combout ),
	.cin(gnd),
	.combout(\reg_file[30][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[30][1]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[30][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N14
cycloneive_lcell_comb \Decoder0~22 (
// Equation(s):
// \Decoder0~22_combout  = (!\prif.regwrite_wb [0] & (\prif.Regwen_wb~q  & \prif.regwrite_wb [2]))

	.dataa(gnd),
	.datab(prifregwrite_wb_0),
	.datac(prifRegwen_wb),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\Decoder0~22_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~22 .lut_mask = 16'h3000;
defparam \Decoder0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N28
cycloneive_lcell_comb \Decoder0~25 (
// Equation(s):
// \Decoder0~25_combout  = (\prif.regwrite_wb [3] & (\prif.regwrite_wb [1] & (\Decoder0~22_combout  & \prif.regwrite_wb [4])))

	.dataa(prifregwrite_wb_3),
	.datab(prifregwrite_wb_1),
	.datac(\Decoder0~22_combout ),
	.datad(prifregwrite_wb_4),
	.cin(gnd),
	.combout(\Decoder0~25_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~25 .lut_mask = 16'h8000;
defparam \Decoder0~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N25
dffeas \reg_file[30][1] (
	.clk(!CLK),
	.d(\reg_file[30][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][1] .is_wysiwyg = "true";
defparam \reg_file[30][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y31_N26
cycloneive_lcell_comb \Decoder0~20 (
// Equation(s):
// \Decoder0~20_combout  = (\prif.Regwen_wb~q  & (!\prif.regwrite_wb [0] & !\prif.regwrite_wb [2]))

	.dataa(prifRegwen_wb),
	.datab(gnd),
	.datac(prifregwrite_wb_0),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\Decoder0~20_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~20 .lut_mask = 16'h000A;
defparam \Decoder0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N22
cycloneive_lcell_comb \Decoder0~24 (
// Equation(s):
// \Decoder0~24_combout  = (\prif.regwrite_wb [1] & (\prif.regwrite_wb [4] & (!\prif.regwrite_wb [3] & \Decoder0~20_combout )))

	.dataa(prifregwrite_wb_1),
	.datab(prifregwrite_wb_4),
	.datac(prifregwrite_wb_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~24_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~24 .lut_mask = 16'h0800;
defparam \Decoder0~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y30_N21
dffeas \reg_file[18][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][1] .is_wysiwyg = "true";
defparam \reg_file[18][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N12
cycloneive_lcell_comb \Decoder0~23 (
// Equation(s):
// \Decoder0~23_combout  = (!\prif.regwrite_wb [3] & (\prif.regwrite_wb [1] & (\Decoder0~22_combout  & \prif.regwrite_wb [4])))

	.dataa(prifregwrite_wb_3),
	.datab(prifregwrite_wb_1),
	.datac(\Decoder0~22_combout ),
	.datad(prifregwrite_wb_4),
	.cin(gnd),
	.combout(\Decoder0~23_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~23 .lut_mask = 16'h4000;
defparam \Decoder0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N29
dffeas \reg_file[22][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][1] .is_wysiwyg = "true";
defparam \reg_file[22][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N20
cycloneive_lcell_comb \Mux62~2 (
// Equation(s):
// \Mux62~2_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[22][1]~q ))) # (!\prif.imemload_id [18] & (\reg_file[18][1]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][1]~q ),
	.datad(\reg_file[22][1]~q ),
	.cin(gnd),
	.combout(\Mux62~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~2 .lut_mask = 16'hDC98;
defparam \Mux62~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N16
cycloneive_lcell_comb \Decoder0~21 (
// Equation(s):
// \Decoder0~21_combout  = (\prif.regwrite_wb [1] & (\prif.regwrite_wb [4] & (\prif.regwrite_wb [3] & \Decoder0~20_combout )))

	.dataa(prifregwrite_wb_1),
	.datab(prifregwrite_wb_4),
	.datac(prifregwrite_wb_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~21_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~21 .lut_mask = 16'h8000;
defparam \Decoder0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N25
dffeas \reg_file[26][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][1] .is_wysiwyg = "true";
defparam \reg_file[26][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N26
cycloneive_lcell_comb \Mux62~3 (
// Equation(s):
// \Mux62~3_combout  = (\prif.imemload_id [19] & ((\Mux62~2_combout  & (\reg_file[30][1]~q )) # (!\Mux62~2_combout  & ((\reg_file[26][1]~q ))))) # (!\prif.imemload_id [19] & (((\Mux62~2_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[30][1]~q ),
	.datac(\Mux62~2_combout ),
	.datad(\reg_file[26][1]~q ),
	.cin(gnd),
	.combout(\Mux62~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~3 .lut_mask = 16'hDAD0;
defparam \Mux62~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N10
cycloneive_lcell_comb \Decoder0~26 (
// Equation(s):
// \Decoder0~26_combout  = (!\prif.regwrite_wb [1] & (\prif.regwrite_wb [4] & (\prif.regwrite_wb [3] & \Decoder0~20_combout )))

	.dataa(prifregwrite_wb_1),
	.datab(prifregwrite_wb_4),
	.datac(prifregwrite_wb_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~26_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~26 .lut_mask = 16'h4000;
defparam \Decoder0~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N5
dffeas \reg_file[24][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][1] .is_wysiwyg = "true";
defparam \reg_file[24][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N20
cycloneive_lcell_comb \Decoder0~27 (
// Equation(s):
// \Decoder0~27_combout  = (!\prif.regwrite_wb [3] & (!\prif.regwrite_wb [1] & (\Decoder0~22_combout  & \prif.regwrite_wb [4])))

	.dataa(prifregwrite_wb_3),
	.datab(prifregwrite_wb_1),
	.datac(\Decoder0~22_combout ),
	.datad(prifregwrite_wb_4),
	.cin(gnd),
	.combout(\Decoder0~27_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~27 .lut_mask = 16'h1000;
defparam \Decoder0~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N13
dffeas \reg_file[20][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][1] .is_wysiwyg = "true";
defparam \reg_file[20][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N18
cycloneive_lcell_comb \Decoder0~28 (
// Equation(s):
// \Decoder0~28_combout  = (!\prif.regwrite_wb [1] & (\prif.regwrite_wb [4] & (!\prif.regwrite_wb [3] & \Decoder0~20_combout )))

	.dataa(prifregwrite_wb_1),
	.datab(prifregwrite_wb_4),
	.datac(prifregwrite_wb_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~28_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~28 .lut_mask = 16'h0400;
defparam \Decoder0~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N3
dffeas \reg_file[16][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][1] .is_wysiwyg = "true";
defparam \reg_file[16][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N12
cycloneive_lcell_comb \Mux62~4 (
// Equation(s):
// \Mux62~4_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[20][1]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[16][1]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[20][1]~q ),
	.datad(\reg_file[16][1]~q ),
	.cin(gnd),
	.combout(\Mux62~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~4 .lut_mask = 16'hB9A8;
defparam \Mux62~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N4
cycloneive_lcell_comb \Mux62~5 (
// Equation(s):
// \Mux62~5_combout  = (\prif.imemload_id [19] & ((\Mux62~4_combout  & (\reg_file[28][1]~q )) # (!\Mux62~4_combout  & ((\reg_file[24][1]~q ))))) # (!\prif.imemload_id [19] & (((\Mux62~4_combout ))))

	.dataa(\reg_file[28][1]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[24][1]~q ),
	.datad(\Mux62~4_combout ),
	.cin(gnd),
	.combout(\Mux62~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~5 .lut_mask = 16'hBBC0;
defparam \Mux62~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N8
cycloneive_lcell_comb \Mux62~6 (
// Equation(s):
// \Mux62~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux62~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & ((\Mux62~5_combout ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux62~3_combout ),
	.datad(\Mux62~5_combout ),
	.cin(gnd),
	.combout(\Mux62~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~6 .lut_mask = 16'hB9A8;
defparam \Mux62~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N20
cycloneive_lcell_comb \reg_file[23][1]~feeder (
// Equation(s):
// \reg_file[23][1]~feeder_combout  = \reg_file_nxt[31][1]~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][1]~64_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[23][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][1]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[23][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N8
cycloneive_lcell_comb \Decoder0~30 (
// Equation(s):
// \Decoder0~30_combout  = (!\prif.regwrite_wb [3] & (\Decoder0~14_combout  & (\prif.regwrite_wb [4] & \prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~14_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~30_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~30 .lut_mask = 16'h4000;
defparam \Decoder0~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N21
dffeas \reg_file[23][1] (
	.clk(!CLK),
	.d(\reg_file[23][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][1] .is_wysiwyg = "true";
defparam \reg_file[23][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N30
cycloneive_lcell_comb \Decoder0~33 (
// Equation(s):
// \Decoder0~33_combout  = (\prif.regwrite_wb [3] & (\Decoder0~14_combout  & (\prif.regwrite_wb [4] & \prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~14_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~33_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~33 .lut_mask = 16'h8000;
defparam \Decoder0~33 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y26_N31
dffeas \reg_file[31][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][1] .is_wysiwyg = "true";
defparam \reg_file[31][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N14
cycloneive_lcell_comb \Decoder0~31 (
// Equation(s):
// \Decoder0~31_combout  = (\prif.regwrite_wb [1] & (\Decoder0~16_combout  & (\prif.regwrite_wb [4] & \prif.regwrite_wb [3])))

	.dataa(prifregwrite_wb_1),
	.datab(\Decoder0~16_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_3),
	.cin(gnd),
	.combout(\Decoder0~31_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~31 .lut_mask = 16'h8000;
defparam \Decoder0~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y26_N25
dffeas \reg_file[27][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][1] .is_wysiwyg = "true";
defparam \reg_file[27][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N16
cycloneive_lcell_comb \Decoder0~32 (
// Equation(s):
// \Decoder0~32_combout  = (\prif.regwrite_wb [1] & (\Decoder0~16_combout  & (\prif.regwrite_wb [4] & !\prif.regwrite_wb [3])))

	.dataa(prifregwrite_wb_1),
	.datab(\Decoder0~16_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_3),
	.cin(gnd),
	.combout(\Decoder0~32_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~32 .lut_mask = 16'h0080;
defparam \Decoder0~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N9
dffeas \reg_file[19][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][1] .is_wysiwyg = "true";
defparam \reg_file[19][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N24
cycloneive_lcell_comb \Mux62~7 (
// Equation(s):
// \Mux62~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][1]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][1]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][1]~q ),
	.datad(\reg_file[19][1]~q ),
	.cin(gnd),
	.combout(\Mux62~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~7 .lut_mask = 16'hD9C8;
defparam \Mux62~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N30
cycloneive_lcell_comb \Mux62~8 (
// Equation(s):
// \Mux62~8_combout  = (\prif.imemload_id [18] & ((\Mux62~7_combout  & ((\reg_file[31][1]~q ))) # (!\Mux62~7_combout  & (\reg_file[23][1]~q )))) # (!\prif.imemload_id [18] & (((\Mux62~7_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[23][1]~q ),
	.datac(\reg_file[31][1]~q ),
	.datad(\Mux62~7_combout ),
	.cin(gnd),
	.combout(\Mux62~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~8 .lut_mask = 16'hF588;
defparam \Mux62~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N6
cycloneive_lcell_comb \Decoder0~47 (
// Equation(s):
// \Decoder0~47_combout  = (!\prif.regwrite_wb [1] & (\Decoder0~16_combout  & (!\prif.regwrite_wb [4] & !\prif.regwrite_wb [3])))

	.dataa(prifregwrite_wb_1),
	.datab(\Decoder0~16_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_3),
	.cin(gnd),
	.combout(\Decoder0~47_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~47 .lut_mask = 16'h0004;
defparam \Decoder0~47 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y27_N19
dffeas \reg_file[1][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][1] .is_wysiwyg = "true";
defparam \reg_file[1][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N12
cycloneive_lcell_comb \reg_file[3][1]~feeder (
// Equation(s):
// \reg_file[3][1]~feeder_combout  = \reg_file_nxt[31][1]~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][1]~64_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[3][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[3][1]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[3][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N24
cycloneive_lcell_comb \Decoder0~46 (
// Equation(s):
// \Decoder0~46_combout  = (\prif.regwrite_wb [1] & (\Decoder0~16_combout  & (!\prif.regwrite_wb [4] & !\prif.regwrite_wb [3])))

	.dataa(prifregwrite_wb_1),
	.datab(\Decoder0~16_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_3),
	.cin(gnd),
	.combout(\Decoder0~46_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~46 .lut_mask = 16'h0008;
defparam \Decoder0~46 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y27_N13
dffeas \reg_file[3][1] (
	.clk(!CLK),
	.d(\reg_file[3][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][1] .is_wysiwyg = "true";
defparam \reg_file[3][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N18
cycloneive_lcell_comb \Mux62~14 (
// Equation(s):
// \Mux62~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][1]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][1]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][1]~q ),
	.datad(\reg_file[3][1]~q ),
	.cin(gnd),
	.combout(\Mux62~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~14 .lut_mask = 16'hC840;
defparam \Mux62~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N2
cycloneive_lcell_comb \Decoder0~48 (
// Equation(s):
// \Decoder0~48_combout  = (\prif.regwrite_wb [1] & (!\prif.regwrite_wb [4] & (!\prif.regwrite_wb [3] & \Decoder0~20_combout )))

	.dataa(prifregwrite_wb_1),
	.datab(prifregwrite_wb_4),
	.datac(prifregwrite_wb_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~48_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~48 .lut_mask = 16'h0200;
defparam \Decoder0~48 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y26_N31
dffeas \reg_file[2][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][1] .is_wysiwyg = "true";
defparam \reg_file[2][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N28
cycloneive_lcell_comb \Mux62~15 (
// Equation(s):
// \Mux62~15_combout  = (\Mux62~14_combout ) # ((\prif.imemload_id [17] & (!\prif.imemload_id [16] & \reg_file[2][1]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux62~14_combout ),
	.datad(\reg_file[2][1]~q ),
	.cin(gnd),
	.combout(\Mux62~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~15 .lut_mask = 16'hF2F0;
defparam \Mux62~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N28
cycloneive_lcell_comb \Decoder0~34 (
// Equation(s):
// \Decoder0~34_combout  = (\prif.regwrite_wb [3] & (\Decoder0~16_combout  & (!\prif.regwrite_wb [4] & !\prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~16_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~34_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~34 .lut_mask = 16'h0008;
defparam \Decoder0~34 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y25_N1
dffeas \reg_file[9][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][1] .is_wysiwyg = "true";
defparam \reg_file[9][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N26
cycloneive_lcell_comb \Decoder0~37 (
// Equation(s):
// \Decoder0~37_combout  = (\Decoder0~16_combout  & (!\prif.regwrite_wb [4] & (\prif.regwrite_wb [3] & \prif.regwrite_wb [1])))

	.dataa(\Decoder0~16_combout ),
	.datab(prifregwrite_wb_4),
	.datac(prifregwrite_wb_3),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~37_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~37 .lut_mask = 16'h2000;
defparam \Decoder0~37 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y25_N23
dffeas \reg_file[11][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][1] .is_wysiwyg = "true";
defparam \reg_file[11][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N6
cycloneive_lcell_comb \Decoder0~35 (
// Equation(s):
// \Decoder0~35_combout  = (\prif.regwrite_wb [1] & (!\prif.regwrite_wb [4] & (\prif.regwrite_wb [3] & \Decoder0~20_combout )))

	.dataa(prifregwrite_wb_1),
	.datab(prifregwrite_wb_4),
	.datac(prifregwrite_wb_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~35_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~35 .lut_mask = 16'h2000;
defparam \Decoder0~35 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y25_N5
dffeas \reg_file[10][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][1] .is_wysiwyg = "true";
defparam \reg_file[10][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N4
cycloneive_lcell_comb \Mux62~12 (
// Equation(s):
// \Mux62~12_combout  = (\prif.imemload_id [17] & (((\reg_file[10][1]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][1]~q  & ((!\prif.imemload_id [16]))))

	.dataa(\reg_file[8][1]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[10][1]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux62~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~12 .lut_mask = 16'hCCE2;
defparam \Mux62~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N22
cycloneive_lcell_comb \Mux62~13 (
// Equation(s):
// \Mux62~13_combout  = (\prif.imemload_id [16] & ((\Mux62~12_combout  & ((\reg_file[11][1]~q ))) # (!\Mux62~12_combout  & (\reg_file[9][1]~q )))) # (!\prif.imemload_id [16] & (((\Mux62~12_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[9][1]~q ),
	.datac(\reg_file[11][1]~q ),
	.datad(\Mux62~12_combout ),
	.cin(gnd),
	.combout(\Mux62~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~13 .lut_mask = 16'hF588;
defparam \Mux62~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N30
cycloneive_lcell_comb \Mux62~16 (
// Equation(s):
// \Mux62~16_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18]) # (\Mux62~13_combout )))) # (!\prif.imemload_id [19] & (\Mux62~15_combout  & (!\prif.imemload_id [18])))

	.dataa(prifimemload_id_19),
	.datab(\Mux62~15_combout ),
	.datac(prifimemload_id_18),
	.datad(\Mux62~13_combout ),
	.cin(gnd),
	.combout(\Mux62~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~16 .lut_mask = 16'hAEA4;
defparam \Mux62~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N10
cycloneive_lcell_comb \Decoder0~39 (
// Equation(s):
// \Decoder0~39_combout  = (\prif.regwrite_wb [3] & (\Decoder0~14_combout  & (!\prif.regwrite_wb [4] & !\prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~14_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~39_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~39 .lut_mask = 16'h0008;
defparam \Decoder0~39 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y25_N9
dffeas \reg_file[13][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][1] .is_wysiwyg = "true";
defparam \reg_file[13][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N24
cycloneive_lcell_comb \Decoder0~40 (
// Equation(s):
// \Decoder0~40_combout  = (!\prif.regwrite_wb [1] & (\prif.regwrite_wb [3] & (\Decoder0~22_combout  & !\prif.regwrite_wb [4])))

	.dataa(prifregwrite_wb_1),
	.datab(prifregwrite_wb_3),
	.datac(\Decoder0~22_combout ),
	.datad(prifregwrite_wb_4),
	.cin(gnd),
	.combout(\Decoder0~40_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~40 .lut_mask = 16'h0040;
defparam \Decoder0~40 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y25_N3
dffeas \reg_file[12][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][1] .is_wysiwyg = "true";
defparam \reg_file[12][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N8
cycloneive_lcell_comb \Mux62~17 (
// Equation(s):
// \Mux62~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & (\reg_file[13][1]~q )) # (!\prif.imemload_id [16] & ((\reg_file[12][1]~q )))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[13][1]~q ),
	.datad(\reg_file[12][1]~q ),
	.cin(gnd),
	.combout(\Mux62~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~17 .lut_mask = 16'hD9C8;
defparam \Mux62~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N20
cycloneive_lcell_comb \Decoder0~38 (
// Equation(s):
// \Decoder0~38_combout  = (\prif.regwrite_wb [3] & (\Decoder0~22_combout  & (!\prif.regwrite_wb [4] & \prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~22_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~38_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~38 .lut_mask = 16'h0800;
defparam \Decoder0~38 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N5
dffeas \reg_file[14][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][1] .is_wysiwyg = "true";
defparam \reg_file[14][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N28
cycloneive_lcell_comb \Decoder0~41 (
// Equation(s):
// \Decoder0~41_combout  = (\prif.regwrite_wb [3] & (\Decoder0~14_combout  & (!\prif.regwrite_wb [4] & \prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~14_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~41_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~41 .lut_mask = 16'h0800;
defparam \Decoder0~41 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N7
dffeas \reg_file[15][1] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][1]~64_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][1] .is_wysiwyg = "true";
defparam \reg_file[15][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N4
cycloneive_lcell_comb \Mux62~18 (
// Equation(s):
// \Mux62~18_combout  = (\prif.imemload_id [17] & ((\Mux62~17_combout  & ((\reg_file[15][1]~q ))) # (!\Mux62~17_combout  & (\reg_file[14][1]~q )))) # (!\prif.imemload_id [17] & (\Mux62~17_combout ))

	.dataa(prifimemload_id_17),
	.datab(\Mux62~17_combout ),
	.datac(\reg_file[14][1]~q ),
	.datad(\reg_file[15][1]~q ),
	.cin(gnd),
	.combout(\Mux62~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~18 .lut_mask = 16'hEC64;
defparam \Mux62~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N24
cycloneive_lcell_comb \reg_file[7][1]~feeder (
// Equation(s):
// \reg_file[7][1]~feeder_combout  = \reg_file_nxt[31][1]~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][1]~64_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[7][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[7][1]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[7][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N26
cycloneive_lcell_comb \Decoder0~45 (
// Equation(s):
// \Decoder0~45_combout  = (!\prif.regwrite_wb [3] & (\Decoder0~14_combout  & (!\prif.regwrite_wb [4] & \prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~14_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~45_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~45 .lut_mask = 16'h0400;
defparam \Decoder0~45 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y26_N25
dffeas \reg_file[7][1] (
	.clk(!CLK),
	.d(\reg_file[7][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][1] .is_wysiwyg = "true";
defparam \reg_file[7][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N14
cycloneive_lcell_comb \Decoder0~42 (
// Equation(s):
// \Decoder0~42_combout  = (!\prif.regwrite_wb [3] & (!\prif.regwrite_wb [4] & (\Decoder0~22_combout  & \prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(prifregwrite_wb_4),
	.datac(\Decoder0~22_combout ),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~42_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~42 .lut_mask = 16'h1000;
defparam \Decoder0~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N29
dffeas \reg_file[6][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][1] .is_wysiwyg = "true";
defparam \reg_file[6][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N0
cycloneive_lcell_comb \Decoder0~44 (
// Equation(s):
// \Decoder0~44_combout  = (!\prif.regwrite_wb [3] & (\Decoder0~22_combout  & (!\prif.regwrite_wb [4] & !\prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~22_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~44_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~44 .lut_mask = 16'h0004;
defparam \Decoder0~44 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N1
dffeas \reg_file[4][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][1] .is_wysiwyg = "true";
defparam \reg_file[4][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N24
cycloneive_lcell_comb \reg_file[5][1]~feeder (
// Equation(s):
// \reg_file[5][1]~feeder_combout  = \reg_file_nxt[31][1]~64_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][1]~64_combout ),
	.cin(gnd),
	.combout(\reg_file[5][1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[5][1]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[5][1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y28_N22
cycloneive_lcell_comb \Decoder0~43 (
// Equation(s):
// \Decoder0~43_combout  = (!\prif.regwrite_wb [3] & (\Decoder0~14_combout  & (!\prif.regwrite_wb [4] & !\prif.regwrite_wb [1])))

	.dataa(prifregwrite_wb_3),
	.datab(\Decoder0~14_combout ),
	.datac(prifregwrite_wb_4),
	.datad(prifregwrite_wb_1),
	.cin(gnd),
	.combout(\Decoder0~43_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~43 .lut_mask = 16'h0004;
defparam \Decoder0~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N25
dffeas \reg_file[5][1] (
	.clk(!CLK),
	.d(\reg_file[5][1]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][1] .is_wysiwyg = "true";
defparam \reg_file[5][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N6
cycloneive_lcell_comb \Mux62~10 (
// Equation(s):
// \Mux62~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][1]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][1]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][1]~q ),
	.datad(\reg_file[5][1]~q ),
	.cin(gnd),
	.combout(\Mux62~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~10 .lut_mask = 16'hBA98;
defparam \Mux62~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N28
cycloneive_lcell_comb \Mux62~11 (
// Equation(s):
// \Mux62~11_combout  = (\prif.imemload_id [17] & ((\Mux62~10_combout  & (\reg_file[7][1]~q )) # (!\Mux62~10_combout  & ((\reg_file[6][1]~q ))))) # (!\prif.imemload_id [17] & (((\Mux62~10_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[7][1]~q ),
	.datac(\reg_file[6][1]~q ),
	.datad(\Mux62~10_combout ),
	.cin(gnd),
	.combout(\Mux62~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux62~11 .lut_mask = 16'hDDA0;
defparam \Mux62~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N16
cycloneive_lcell_comb \Mux30~0 (
// Equation(s):
// \Mux30~0_combout  = (\prif.imemload_id [23] & (((\reg_file[21][1]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[17][1]~q  & ((!\prif.imemload_id [24]))))

	.dataa(\reg_file[17][1]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[21][1]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux30~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~0 .lut_mask = 16'hCCE2;
defparam \Mux30~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N12
cycloneive_lcell_comb \Mux30~1 (
// Equation(s):
// \Mux30~1_combout  = (\prif.imemload_id [24] & ((\Mux30~0_combout  & (\reg_file[29][1]~q )) # (!\Mux30~0_combout  & ((\reg_file[25][1]~q ))))) # (!\prif.imemload_id [24] & (((\Mux30~0_combout ))))

	.dataa(\reg_file[29][1]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[25][1]~q ),
	.datad(\Mux30~0_combout ),
	.cin(gnd),
	.combout(\Mux30~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~1 .lut_mask = 16'hBBC0;
defparam \Mux30~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N8
cycloneive_lcell_comb \Mux30~7 (
// Equation(s):
// \Mux30~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][1]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][1]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][1]~q ),
	.datad(\reg_file[23][1]~q ),
	.cin(gnd),
	.combout(\Mux30~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~7 .lut_mask = 16'hDC98;
defparam \Mux30~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N30
cycloneive_lcell_comb \Mux30~8 (
// Equation(s):
// \Mux30~8_combout  = (\Mux30~7_combout  & (((\reg_file[31][1]~q ) # (!\prif.imemload_id [24])))) # (!\Mux30~7_combout  & (\reg_file[27][1]~q  & ((\prif.imemload_id [24]))))

	.dataa(\Mux30~7_combout ),
	.datab(\reg_file[27][1]~q ),
	.datac(\reg_file[31][1]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux30~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~8 .lut_mask = 16'hE4AA;
defparam \Mux30~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N24
cycloneive_lcell_comb \Mux30~2 (
// Equation(s):
// \Mux30~2_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[26][1]~q ))) # (!\prif.imemload_id [24] & (\reg_file[18][1]~q ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[18][1]~q ),
	.datac(\reg_file[26][1]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux30~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~2 .lut_mask = 16'hFA44;
defparam \Mux30~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N28
cycloneive_lcell_comb \Mux30~3 (
// Equation(s):
// \Mux30~3_combout  = (\prif.imemload_id [23] & ((\Mux30~2_combout  & (\reg_file[30][1]~q )) # (!\Mux30~2_combout  & ((\reg_file[22][1]~q ))))) # (!\prif.imemload_id [23] & (((\Mux30~2_combout ))))

	.dataa(\reg_file[30][1]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[22][1]~q ),
	.datad(\Mux30~2_combout ),
	.cin(gnd),
	.combout(\Mux30~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~3 .lut_mask = 16'hBBC0;
defparam \Mux30~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N0
cycloneive_lcell_comb \Decoder0~29 (
// Equation(s):
// \Decoder0~29_combout  = (\prif.regwrite_wb [3] & (!\prif.regwrite_wb [1] & (\Decoder0~22_combout  & \prif.regwrite_wb [4])))

	.dataa(prifregwrite_wb_3),
	.datab(prifregwrite_wb_1),
	.datac(\Decoder0~22_combout ),
	.datad(prifregwrite_wb_4),
	.cin(gnd),
	.combout(\Decoder0~29_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~29 .lut_mask = 16'h2000;
defparam \Decoder0~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N31
dffeas \reg_file[28][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][1] .is_wysiwyg = "true";
defparam \reg_file[28][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N30
cycloneive_lcell_comb \Mux30~5 (
// Equation(s):
// \Mux30~5_combout  = (\Mux30~4_combout  & (((\reg_file[28][1]~q )) # (!\prif.imemload_id [23]))) # (!\Mux30~4_combout  & (\prif.imemload_id [23] & ((\reg_file[20][1]~q ))))

	.dataa(\Mux30~4_combout ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[28][1]~q ),
	.datad(\reg_file[20][1]~q ),
	.cin(gnd),
	.combout(\Mux30~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~5 .lut_mask = 16'hE6A2;
defparam \Mux30~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N24
cycloneive_lcell_comb \Mux30~6 (
// Equation(s):
// \Mux30~6_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\Mux30~3_combout )) # (!\prif.imemload_id [22] & ((\Mux30~5_combout )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux30~3_combout ),
	.datad(\Mux30~5_combout ),
	.cin(gnd),
	.combout(\Mux30~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~6 .lut_mask = 16'hD9C8;
defparam \Mux30~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N30
cycloneive_lcell_comb \Mux30~15 (
// Equation(s):
// \Mux30~15_combout  = (\Mux30~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][1]~q  & !\prif.imemload_id [21])))

	.dataa(\Mux30~14_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][1]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux30~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~15 .lut_mask = 16'hAAEA;
defparam \Mux30~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N0
cycloneive_lcell_comb \Mux30~12 (
// Equation(s):
// \Mux30~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][1]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[4][1]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[4][1]~q ),
	.datad(\reg_file[5][1]~q ),
	.cin(gnd),
	.combout(\Mux30~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~12 .lut_mask = 16'hBA98;
defparam \Mux30~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N4
cycloneive_lcell_comb \Mux30~13 (
// Equation(s):
// \Mux30~13_combout  = (\prif.imemload_id [22] & ((\Mux30~12_combout  & (\reg_file[7][1]~q )) # (!\Mux30~12_combout  & ((\reg_file[6][1]~q ))))) # (!\prif.imemload_id [22] & (((\Mux30~12_combout ))))

	.dataa(\reg_file[7][1]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[6][1]~q ),
	.datad(\Mux30~12_combout ),
	.cin(gnd),
	.combout(\Mux30~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~13 .lut_mask = 16'hBBC0;
defparam \Mux30~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N10
cycloneive_lcell_comb \Mux30~16 (
// Equation(s):
// \Mux30~16_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\Mux30~13_combout ))) # (!\prif.imemload_id [23] & (\Mux30~15_combout ))))

	.dataa(\Mux30~15_combout ),
	.datab(prifimemload_id_24),
	.datac(prifimemload_id_23),
	.datad(\Mux30~13_combout ),
	.cin(gnd),
	.combout(\Mux30~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~16 .lut_mask = 16'hF2C2;
defparam \Mux30~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N4
cycloneive_lcell_comb \Decoder0~36 (
// Equation(s):
// \Decoder0~36_combout  = (!\prif.regwrite_wb [1] & (!\prif.regwrite_wb [4] & (\prif.regwrite_wb [3] & \Decoder0~20_combout )))

	.dataa(prifregwrite_wb_1),
	.datab(prifregwrite_wb_4),
	.datac(prifregwrite_wb_3),
	.datad(\Decoder0~20_combout ),
	.cin(gnd),
	.combout(\Decoder0~36_combout ),
	.cout());
// synopsys translate_off
defparam \Decoder0~36 .lut_mask = 16'h1000;
defparam \Decoder0~36 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y25_N23
dffeas \reg_file[8][1] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][1]~64_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][1]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][1] .is_wysiwyg = "true";
defparam \reg_file[8][1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N22
cycloneive_lcell_comb \Mux30~10 (
// Equation(s):
// \Mux30~10_combout  = (\prif.imemload_id [22] & ((\reg_file[10][1]~q ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\reg_file[8][1]~q  & !\prif.imemload_id [21]))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[10][1]~q ),
	.datac(\reg_file[8][1]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux30~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~10 .lut_mask = 16'hAAD8;
defparam \Mux30~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N0
cycloneive_lcell_comb \Mux30~11 (
// Equation(s):
// \Mux30~11_combout  = (\prif.imemload_id [21] & ((\Mux30~10_combout  & (\reg_file[11][1]~q )) # (!\Mux30~10_combout  & ((\reg_file[9][1]~q ))))) # (!\prif.imemload_id [21] & (((\Mux30~10_combout ))))

	.dataa(\reg_file[11][1]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[9][1]~q ),
	.datad(\Mux30~10_combout ),
	.cin(gnd),
	.combout(\Mux30~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~11 .lut_mask = 16'hBBC0;
defparam \Mux30~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N2
cycloneive_lcell_comb \Mux30~17 (
// Equation(s):
// \Mux30~17_combout  = (\prif.imemload_id [21] & ((\reg_file[13][1]~q ) # ((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (((\reg_file[12][1]~q  & !\prif.imemload_id [22]))))

	.dataa(\reg_file[13][1]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[12][1]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux30~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~17 .lut_mask = 16'hCCB8;
defparam \Mux30~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N28
cycloneive_lcell_comb \Mux30~18 (
// Equation(s):
// \Mux30~18_combout  = (\prif.imemload_id [22] & ((\Mux30~17_combout  & (\reg_file[15][1]~q )) # (!\Mux30~17_combout  & ((\reg_file[14][1]~q ))))) # (!\prif.imemload_id [22] & (((\Mux30~17_combout ))))

	.dataa(\reg_file[15][1]~q ),
	.datab(\reg_file[14][1]~q ),
	.datac(prifimemload_id_22),
	.datad(\Mux30~17_combout ),
	.cin(gnd),
	.combout(\Mux30~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux30~18 .lut_mask = 16'hAFC0;
defparam \Mux30~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N24
cycloneive_lcell_comb \reg_file_nxt[31][0]~65 (
// Equation(s):
// \reg_file_nxt[31][0]~65_combout  = (\Mux164~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Mux164),
	.datac(prifregwrite_wb_0),
	.datad(Equal8),
	.cin(gnd),
	.combout(\reg_file_nxt[31][0]~65_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][0]~65 .lut_mask = 16'hC8CC;
defparam \reg_file_nxt[31][0]~65 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N5
dffeas \reg_file[31][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][0] .is_wysiwyg = "true";
defparam \reg_file[31][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N11
dffeas \reg_file[19][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][0] .is_wysiwyg = "true";
defparam \reg_file[19][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N19
dffeas \reg_file[23][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][0] .is_wysiwyg = "true";
defparam \reg_file[23][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N18
cycloneive_lcell_comb \Mux63~7 (
// Equation(s):
// \Mux63~7_combout  = (\prif.imemload_id [18] & (((\reg_file[23][0]~q ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\reg_file[19][0]~q  & ((!\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[19][0]~q ),
	.datac(\reg_file[23][0]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux63~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~7 .lut_mask = 16'hAAE4;
defparam \Mux63~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N25
dffeas \reg_file[27][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][0] .is_wysiwyg = "true";
defparam \reg_file[27][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N24
cycloneive_lcell_comb \Mux63~8 (
// Equation(s):
// \Mux63~8_combout  = (\Mux63~7_combout  & ((\reg_file[31][0]~q ) # ((!\prif.imemload_id [19])))) # (!\Mux63~7_combout  & (((\reg_file[27][0]~q  & \prif.imemload_id [19]))))

	.dataa(\reg_file[31][0]~q ),
	.datab(\Mux63~7_combout ),
	.datac(\reg_file[27][0]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux63~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~8 .lut_mask = 16'hB8CC;
defparam \Mux63~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N24
cycloneive_lcell_comb \reg_file[25][0]~feeder (
// Equation(s):
// \reg_file[25][0]~feeder_combout  = \reg_file_nxt[31][0]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][0]~65_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[25][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][0]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[25][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N25
dffeas \reg_file[25][0] (
	.clk(!CLK),
	.d(\reg_file[25][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][0] .is_wysiwyg = "true";
defparam \reg_file[25][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y31_N25
dffeas \reg_file[29][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][0] .is_wysiwyg = "true";
defparam \reg_file[29][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N31
dffeas \reg_file[17][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][0] .is_wysiwyg = "true";
defparam \reg_file[17][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N24
cycloneive_lcell_comb \reg_file[21][0]~feeder (
// Equation(s):
// \reg_file[21][0]~feeder_combout  = \reg_file_nxt[31][0]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][0]~65_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[21][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][0]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[21][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N25
dffeas \reg_file[21][0] (
	.clk(!CLK),
	.d(\reg_file[21][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][0] .is_wysiwyg = "true";
defparam \reg_file[21][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N26
cycloneive_lcell_comb \Mux63~0 (
// Equation(s):
// \Mux63~0_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19]) # (\reg_file[21][0]~q )))) # (!\prif.imemload_id [18] & (\reg_file[17][0]~q  & (!\prif.imemload_id [19])))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[17][0]~q ),
	.datac(prifimemload_id_19),
	.datad(\reg_file[21][0]~q ),
	.cin(gnd),
	.combout(\Mux63~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~0 .lut_mask = 16'hAEA4;
defparam \Mux63~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N30
cycloneive_lcell_comb \Mux63~1 (
// Equation(s):
// \Mux63~1_combout  = (\prif.imemload_id [19] & ((\Mux63~0_combout  & ((\reg_file[29][0]~q ))) # (!\Mux63~0_combout  & (\reg_file[25][0]~q )))) # (!\prif.imemload_id [19] & (((\Mux63~0_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[25][0]~q ),
	.datac(\reg_file[29][0]~q ),
	.datad(\Mux63~0_combout ),
	.cin(gnd),
	.combout(\Mux63~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~1 .lut_mask = 16'hF588;
defparam \Mux63~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N25
dffeas \reg_file[20][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][0] .is_wysiwyg = "true";
defparam \reg_file[20][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N27
dffeas \reg_file[28][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][0] .is_wysiwyg = "true";
defparam \reg_file[28][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N5
dffeas \reg_file[16][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][0] .is_wysiwyg = "true";
defparam \reg_file[16][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N22
cycloneive_lcell_comb \reg_file[24][0]~feeder (
// Equation(s):
// \reg_file[24][0]~feeder_combout  = \reg_file_nxt[31][0]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][0]~65_combout ),
	.cin(gnd),
	.combout(\reg_file[24][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][0]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[24][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N23
dffeas \reg_file[24][0] (
	.clk(!CLK),
	.d(\reg_file[24][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][0] .is_wysiwyg = "true";
defparam \reg_file[24][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N4
cycloneive_lcell_comb \Mux63~4 (
// Equation(s):
// \Mux63~4_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[24][0]~q ))) # (!\prif.imemload_id [19] & (\reg_file[16][0]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[16][0]~q ),
	.datad(\reg_file[24][0]~q ),
	.cin(gnd),
	.combout(\Mux63~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~4 .lut_mask = 16'hDC98;
defparam \Mux63~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N16
cycloneive_lcell_comb \Mux63~5 (
// Equation(s):
// \Mux63~5_combout  = (\prif.imemload_id [18] & ((\Mux63~4_combout  & ((\reg_file[28][0]~q ))) # (!\Mux63~4_combout  & (\reg_file[20][0]~q )))) # (!\prif.imemload_id [18] & (((\Mux63~4_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[20][0]~q ),
	.datac(\reg_file[28][0]~q ),
	.datad(\Mux63~4_combout ),
	.cin(gnd),
	.combout(\Mux63~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~5 .lut_mask = 16'hF588;
defparam \Mux63~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N9
dffeas \reg_file[22][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][0] .is_wysiwyg = "true";
defparam \reg_file[22][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N11
dffeas \reg_file[18][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][0] .is_wysiwyg = "true";
defparam \reg_file[18][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N0
cycloneive_lcell_comb \reg_file[26][0]~feeder (
// Equation(s):
// \reg_file[26][0]~feeder_combout  = \reg_file_nxt[31][0]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][0]~65_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[26][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[26][0]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[26][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N1
dffeas \reg_file[26][0] (
	.clk(!CLK),
	.d(\reg_file[26][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][0] .is_wysiwyg = "true";
defparam \reg_file[26][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N10
cycloneive_lcell_comb \Mux63~2 (
// Equation(s):
// \Mux63~2_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[26][0]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & (\reg_file[18][0]~q )))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][0]~q ),
	.datad(\reg_file[26][0]~q ),
	.cin(gnd),
	.combout(\Mux63~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~2 .lut_mask = 16'hBA98;
defparam \Mux63~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N8
cycloneive_lcell_comb \Mux63~3 (
// Equation(s):
// \Mux63~3_combout  = (\prif.imemload_id [18] & ((\Mux63~2_combout  & (\reg_file[30][0]~q )) # (!\Mux63~2_combout  & ((\reg_file[22][0]~q ))))) # (!\prif.imemload_id [18] & (((\Mux63~2_combout ))))

	.dataa(\reg_file[30][0]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[22][0]~q ),
	.datad(\Mux63~2_combout ),
	.cin(gnd),
	.combout(\Mux63~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~3 .lut_mask = 16'hBBC0;
defparam \Mux63~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y27_N10
cycloneive_lcell_comb \Mux63~6 (
// Equation(s):
// \Mux63~6_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\Mux63~3_combout ))) # (!\prif.imemload_id [17] & (\Mux63~5_combout ))))

	.dataa(\Mux63~5_combout ),
	.datab(prifimemload_id_16),
	.datac(prifimemload_id_17),
	.datad(\Mux63~3_combout ),
	.cin(gnd),
	.combout(\Mux63~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~6 .lut_mask = 16'hF2C2;
defparam \Mux63~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N17
dffeas \reg_file[14][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][0] .is_wysiwyg = "true";
defparam \reg_file[14][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N1
dffeas \reg_file[13][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][0] .is_wysiwyg = "true";
defparam \reg_file[13][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N7
dffeas \reg_file[12][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][0] .is_wysiwyg = "true";
defparam \reg_file[12][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N0
cycloneive_lcell_comb \Mux63~17 (
// Equation(s):
// \Mux63~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & (\reg_file[13][0]~q )) # (!\prif.imemload_id [16] & ((\reg_file[12][0]~q )))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[13][0]~q ),
	.datad(\reg_file[12][0]~q ),
	.cin(gnd),
	.combout(\Mux63~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~17 .lut_mask = 16'hD9C8;
defparam \Mux63~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N25
dffeas \reg_file[15][0] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][0]~65_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][0] .is_wysiwyg = "true";
defparam \reg_file[15][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N12
cycloneive_lcell_comb \Mux63~18 (
// Equation(s):
// \Mux63~18_combout  = (\prif.imemload_id [17] & ((\Mux63~17_combout  & ((\reg_file[15][0]~q ))) # (!\Mux63~17_combout  & (\reg_file[14][0]~q )))) # (!\prif.imemload_id [17] & (((\Mux63~17_combout ))))

	.dataa(\reg_file[14][0]~q ),
	.datab(prifimemload_id_17),
	.datac(\Mux63~17_combout ),
	.datad(\reg_file[15][0]~q ),
	.cin(gnd),
	.combout(\Mux63~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~18 .lut_mask = 16'hF838;
defparam \Mux63~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N0
cycloneive_lcell_comb \reg_file[6][0]~feeder (
// Equation(s):
// \reg_file[6][0]~feeder_combout  = \reg_file_nxt[31][0]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][0]~65_combout ),
	.cin(gnd),
	.combout(\reg_file[6][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][0]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[6][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N1
dffeas \reg_file[6][0] (
	.clk(!CLK),
	.d(\reg_file[6][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][0] .is_wysiwyg = "true";
defparam \reg_file[6][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N16
cycloneive_lcell_comb \reg_file[7][0]~feeder (
// Equation(s):
// \reg_file[7][0]~feeder_combout  = \reg_file_nxt[31][0]~65_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][0]~65_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[7][0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[7][0]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[7][0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y27_N17
dffeas \reg_file[7][0] (
	.clk(!CLK),
	.d(\reg_file[7][0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][0] .is_wysiwyg = "true";
defparam \reg_file[7][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N22
cycloneive_lcell_comb \Mux63~13 (
// Equation(s):
// \Mux63~13_combout  = (\Mux63~12_combout  & (((\reg_file[7][0]~q )) # (!\prif.imemload_id [17]))) # (!\Mux63~12_combout  & (\prif.imemload_id [17] & (\reg_file[6][0]~q )))

	.dataa(\Mux63~12_combout ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[6][0]~q ),
	.datad(\reg_file[7][0]~q ),
	.cin(gnd),
	.combout(\Mux63~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~13 .lut_mask = 16'hEA62;
defparam \Mux63~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y27_N21
dffeas \reg_file[2][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][0] .is_wysiwyg = "true";
defparam \reg_file[2][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y25_N9
dffeas \reg_file[3][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][0] .is_wysiwyg = "true";
defparam \reg_file[3][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y25_N15
dffeas \reg_file[1][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][0] .is_wysiwyg = "true";
defparam \reg_file[1][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N14
cycloneive_lcell_comb \Mux63~14 (
// Equation(s):
// \Mux63~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][0]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][0]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[3][0]~q ),
	.datac(\reg_file[1][0]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux63~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~14 .lut_mask = 16'hD800;
defparam \Mux63~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N20
cycloneive_lcell_comb \Mux63~15 (
// Equation(s):
// \Mux63~15_combout  = (\Mux63~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][0]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[2][0]~q ),
	.datad(\Mux63~14_combout ),
	.cin(gnd),
	.combout(\Mux63~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~15 .lut_mask = 16'hFF40;
defparam \Mux63~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N14
cycloneive_lcell_comb \Mux63~16 (
// Equation(s):
// \Mux63~16_combout  = (\prif.imemload_id [18] & ((\Mux63~13_combout ) # ((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (((\Mux63~15_combout  & !\prif.imemload_id [19]))))

	.dataa(\Mux63~13_combout ),
	.datab(\Mux63~15_combout ),
	.datac(prifimemload_id_18),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux63~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~16 .lut_mask = 16'hF0AC;
defparam \Mux63~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y25_N15
dffeas \reg_file[11][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][0] .is_wysiwyg = "true";
defparam \reg_file[11][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y25_N9
dffeas \reg_file[9][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][0] .is_wysiwyg = "true";
defparam \reg_file[9][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N13
dffeas \reg_file[10][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][0] .is_wysiwyg = "true";
defparam \reg_file[10][0] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N3
dffeas \reg_file[8][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][0] .is_wysiwyg = "true";
defparam \reg_file[8][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N12
cycloneive_lcell_comb \Mux63~10 (
// Equation(s):
// \Mux63~10_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[10][0]~q )) # (!\prif.imemload_id [17] & ((\reg_file[8][0]~q )))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[10][0]~q ),
	.datad(\reg_file[8][0]~q ),
	.cin(gnd),
	.combout(\Mux63~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~10 .lut_mask = 16'hD9C8;
defparam \Mux63~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N8
cycloneive_lcell_comb \Mux63~11 (
// Equation(s):
// \Mux63~11_combout  = (\prif.imemload_id [16] & ((\Mux63~10_combout  & (\reg_file[11][0]~q )) # (!\Mux63~10_combout  & ((\reg_file[9][0]~q ))))) # (!\prif.imemload_id [16] & (((\Mux63~10_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[11][0]~q ),
	.datac(\reg_file[9][0]~q ),
	.datad(\Mux63~10_combout ),
	.cin(gnd),
	.combout(\Mux63~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux63~11 .lut_mask = 16'hDDA0;
defparam \Mux63~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N10
cycloneive_lcell_comb \Mux31~7 (
// Equation(s):
// \Mux31~7_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[27][0]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[19][0]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][0]~q ),
	.datad(\reg_file[27][0]~q ),
	.cin(gnd),
	.combout(\Mux31~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~7 .lut_mask = 16'hBA98;
defparam \Mux31~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N4
cycloneive_lcell_comb \Mux31~8 (
// Equation(s):
// \Mux31~8_combout  = (\Mux31~7_combout  & (((\reg_file[31][0]~q )) # (!\prif.imemload_id [23]))) # (!\Mux31~7_combout  & (\prif.imemload_id [23] & ((\reg_file[23][0]~q ))))

	.dataa(\Mux31~7_combout ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[31][0]~q ),
	.datad(\reg_file[23][0]~q ),
	.cin(gnd),
	.combout(\Mux31~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~8 .lut_mask = 16'hE6A2;
defparam \Mux31~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N24
cycloneive_lcell_comb \Mux31~4 (
// Equation(s):
// \Mux31~4_combout  = (\prif.imemload_id [23] & (((\reg_file[20][0]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[16][0]~q  & ((!\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[16][0]~q ),
	.datac(\reg_file[20][0]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux31~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~4 .lut_mask = 16'hAAE4;
defparam \Mux31~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N26
cycloneive_lcell_comb \Mux31~5 (
// Equation(s):
// \Mux31~5_combout  = (\prif.imemload_id [24] & ((\Mux31~4_combout  & ((\reg_file[28][0]~q ))) # (!\Mux31~4_combout  & (\reg_file[24][0]~q )))) # (!\prif.imemload_id [24] & (((\Mux31~4_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[24][0]~q ),
	.datac(\reg_file[28][0]~q ),
	.datad(\Mux31~4_combout ),
	.cin(gnd),
	.combout(\Mux31~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~5 .lut_mask = 16'hF588;
defparam \Mux31~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N8
cycloneive_lcell_comb \Mux31~2 (
// Equation(s):
// \Mux31~2_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\reg_file[22][0]~q )) # (!\prif.imemload_id [23] & ((\reg_file[18][0]~q )))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[22][0]~q ),
	.datad(\reg_file[18][0]~q ),
	.cin(gnd),
	.combout(\Mux31~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~2 .lut_mask = 16'hD9C8;
defparam \Mux31~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N17
dffeas \reg_file[30][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][0] .is_wysiwyg = "true";
defparam \reg_file[30][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N16
cycloneive_lcell_comb \Mux31~3 (
// Equation(s):
// \Mux31~3_combout  = (\prif.imemload_id [24] & ((\Mux31~2_combout  & (\reg_file[30][0]~q )) # (!\Mux31~2_combout  & ((\reg_file[26][0]~q ))))) # (!\prif.imemload_id [24] & (\Mux31~2_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux31~2_combout ),
	.datac(\reg_file[30][0]~q ),
	.datad(\reg_file[26][0]~q ),
	.cin(gnd),
	.combout(\Mux31~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~3 .lut_mask = 16'hE6C4;
defparam \Mux31~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N24
cycloneive_lcell_comb \Mux31~6 (
// Equation(s):
// \Mux31~6_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21]) # (\Mux31~3_combout )))) # (!\prif.imemload_id [22] & (\Mux31~5_combout  & (!\prif.imemload_id [21])))

	.dataa(prifimemload_id_22),
	.datab(\Mux31~5_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux31~3_combout ),
	.cin(gnd),
	.combout(\Mux31~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~6 .lut_mask = 16'hAEA4;
defparam \Mux31~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N30
cycloneive_lcell_comb \Mux31~0 (
// Equation(s):
// \Mux31~0_combout  = (\prif.imemload_id [24] & ((\reg_file[25][0]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[17][0]~q  & !\prif.imemload_id [23]))))

	.dataa(\reg_file[25][0]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[17][0]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux31~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~0 .lut_mask = 16'hCCB8;
defparam \Mux31~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N24
cycloneive_lcell_comb \Mux31~1 (
// Equation(s):
// \Mux31~1_combout  = (\prif.imemload_id [23] & ((\Mux31~0_combout  & (\reg_file[29][0]~q )) # (!\Mux31~0_combout  & ((\reg_file[21][0]~q ))))) # (!\prif.imemload_id [23] & (\Mux31~0_combout ))

	.dataa(prifimemload_id_23),
	.datab(\Mux31~0_combout ),
	.datac(\reg_file[29][0]~q ),
	.datad(\reg_file[21][0]~q ),
	.cin(gnd),
	.combout(\Mux31~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~1 .lut_mask = 16'hE6C4;
defparam \Mux31~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N14
cycloneive_lcell_comb \Mux31~13 (
// Equation(s):
// \Mux31~13_combout  = (\Mux31~12_combout  & (((\reg_file[11][0]~q ) # (!\prif.imemload_id [21])))) # (!\Mux31~12_combout  & (\reg_file[9][0]~q  & ((\prif.imemload_id [21]))))

	.dataa(\Mux31~12_combout ),
	.datab(\reg_file[9][0]~q ),
	.datac(\reg_file[11][0]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux31~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~13 .lut_mask = 16'hE4AA;
defparam \Mux31~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N8
cycloneive_lcell_comb \Mux31~14 (
// Equation(s):
// \Mux31~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][0]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][0]~q ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[1][0]~q ),
	.datac(\reg_file[3][0]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux31~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~14 .lut_mask = 16'hA088;
defparam \Mux31~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N16
cycloneive_lcell_comb \Mux31~15 (
// Equation(s):
// \Mux31~15_combout  = (\Mux31~14_combout ) # ((!\prif.imemload_id [21] & (\prif.imemload_id [22] & \reg_file[2][0]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux31~14_combout ),
	.datad(\reg_file[2][0]~q ),
	.cin(gnd),
	.combout(\Mux31~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~15 .lut_mask = 16'hF4F0;
defparam \Mux31~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N18
cycloneive_lcell_comb \Mux31~16 (
// Equation(s):
// \Mux31~16_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\Mux31~13_combout )) # (!\prif.imemload_id [24] & ((\Mux31~15_combout )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux31~13_combout ),
	.datad(\Mux31~15_combout ),
	.cin(gnd),
	.combout(\Mux31~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~16 .lut_mask = 16'hD9C8;
defparam \Mux31~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N6
cycloneive_lcell_comb \Mux31~17 (
// Equation(s):
// \Mux31~17_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[13][0]~q ))) # (!\prif.imemload_id [21] & (\reg_file[12][0]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[12][0]~q ),
	.datad(\reg_file[13][0]~q ),
	.cin(gnd),
	.combout(\Mux31~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~17 .lut_mask = 16'hDC98;
defparam \Mux31~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N16
cycloneive_lcell_comb \Mux31~18 (
// Equation(s):
// \Mux31~18_combout  = (\prif.imemload_id [22] & ((\Mux31~17_combout  & (\reg_file[15][0]~q )) # (!\Mux31~17_combout  & ((\reg_file[14][0]~q ))))) # (!\prif.imemload_id [22] & (((\Mux31~17_combout ))))

	.dataa(\reg_file[15][0]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[14][0]~q ),
	.datad(\Mux31~17_combout ),
	.cin(gnd),
	.combout(\Mux31~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~18 .lut_mask = 16'hBBC0;
defparam \Mux31~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y26_N1
dffeas \reg_file[5][0] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][0]~65_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][0]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][0] .is_wysiwyg = "true";
defparam \reg_file[5][0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N0
cycloneive_lcell_comb \Mux31~10 (
// Equation(s):
// \Mux31~10_combout  = (\prif.imemload_id [21] & (((\reg_file[5][0]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[4][0]~q  & ((!\prif.imemload_id [22]))))

	.dataa(\reg_file[4][0]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[5][0]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux31~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~10 .lut_mask = 16'hCCE2;
defparam \Mux31~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N10
cycloneive_lcell_comb \Mux31~11 (
// Equation(s):
// \Mux31~11_combout  = (\prif.imemload_id [22] & ((\Mux31~10_combout  & (\reg_file[7][0]~q )) # (!\Mux31~10_combout  & ((\reg_file[6][0]~q ))))) # (!\prif.imemload_id [22] & (((\Mux31~10_combout ))))

	.dataa(\reg_file[7][0]~q ),
	.datab(\reg_file[6][0]~q ),
	.datac(prifimemload_id_22),
	.datad(\Mux31~10_combout ),
	.cin(gnd),
	.combout(\Mux31~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux31~11 .lut_mask = 16'hAFC0;
defparam \Mux31~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N28
cycloneive_lcell_comb \reg_file_nxt[31][3]~66 (
// Equation(s):
// \reg_file_nxt[31][3]~66_combout  = (\Mux161~1_combout  & ((\prif.regwrite_wb [0]) # ((\prif.regwrite_wb [2]) # (!Equal8))))

	.dataa(Mux161),
	.datab(prifregwrite_wb_0),
	.datac(Equal8),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\reg_file_nxt[31][3]~66_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][3]~66 .lut_mask = 16'hAA8A;
defparam \reg_file_nxt[31][3]~66 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y26_N27
dffeas \reg_file[31][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][3] .is_wysiwyg = "true";
defparam \reg_file[31][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N13
dffeas \reg_file[23][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][3] .is_wysiwyg = "true";
defparam \reg_file[23][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y26_N1
dffeas \reg_file[27][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][3] .is_wysiwyg = "true";
defparam \reg_file[27][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N31
dffeas \reg_file[19][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][3] .is_wysiwyg = "true";
defparam \reg_file[19][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N0
cycloneive_lcell_comb \Mux60~7 (
// Equation(s):
// \Mux60~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][3]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][3]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][3]~q ),
	.datad(\reg_file[19][3]~q ),
	.cin(gnd),
	.combout(\Mux60~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~7 .lut_mask = 16'hD9C8;
defparam \Mux60~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N12
cycloneive_lcell_comb \Mux60~8 (
// Equation(s):
// \Mux60~8_combout  = (\prif.imemload_id [18] & ((\Mux60~7_combout  & (\reg_file[31][3]~q )) # (!\Mux60~7_combout  & ((\reg_file[23][3]~q ))))) # (!\prif.imemload_id [18] & (((\Mux60~7_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[31][3]~q ),
	.datac(\reg_file[23][3]~q ),
	.datad(\Mux60~7_combout ),
	.cin(gnd),
	.combout(\Mux60~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~8 .lut_mask = 16'hDDA0;
defparam \Mux60~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N24
cycloneive_lcell_comb \reg_file[29][3]~feeder (
// Equation(s):
// \reg_file[29][3]~feeder_combout  = \reg_file_nxt[31][3]~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][3]~66_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][3]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N25
dffeas \reg_file[29][3] (
	.clk(!CLK),
	.d(\reg_file[29][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][3] .is_wysiwyg = "true";
defparam \reg_file[29][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N3
dffeas \reg_file[21][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][3] .is_wysiwyg = "true";
defparam \reg_file[21][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N26
cycloneive_lcell_comb \reg_file[25][3]~feeder (
// Equation(s):
// \reg_file[25][3]~feeder_combout  = \reg_file_nxt[31][3]~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][3]~66_combout ),
	.cin(gnd),
	.combout(\reg_file[25][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][3]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[25][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N27
dffeas \reg_file[25][3] (
	.clk(!CLK),
	.d(\reg_file[25][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][3] .is_wysiwyg = "true";
defparam \reg_file[25][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N26
cycloneive_lcell_comb \reg_file[17][3]~feeder (
// Equation(s):
// \reg_file[17][3]~feeder_combout  = \reg_file_nxt[31][3]~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][3]~66_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[17][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[17][3]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[17][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N27
dffeas \reg_file[17][3] (
	.clk(!CLK),
	.d(\reg_file[17][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][3] .is_wysiwyg = "true";
defparam \reg_file[17][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N24
cycloneive_lcell_comb \Mux60~0 (
// Equation(s):
// \Mux60~0_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[25][3]~q )) # (!\prif.imemload_id [19] & ((\reg_file[17][3]~q )))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[25][3]~q ),
	.datac(\reg_file[17][3]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux60~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~0 .lut_mask = 16'hEE50;
defparam \Mux60~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N2
cycloneive_lcell_comb \Mux60~1 (
// Equation(s):
// \Mux60~1_combout  = (\prif.imemload_id [18] & ((\Mux60~0_combout  & (\reg_file[29][3]~q )) # (!\Mux60~0_combout  & ((\reg_file[21][3]~q ))))) # (!\prif.imemload_id [18] & (((\Mux60~0_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[29][3]~q ),
	.datac(\reg_file[21][3]~q ),
	.datad(\Mux60~0_combout ),
	.cin(gnd),
	.combout(\Mux60~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~1 .lut_mask = 16'hDDA0;
defparam \Mux60~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N4
cycloneive_lcell_comb \reg_file[30][3]~feeder (
// Equation(s):
// \reg_file[30][3]~feeder_combout  = \reg_file_nxt[31][3]~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][3]~66_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[30][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[30][3]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[30][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y30_N5
dffeas \reg_file[30][3] (
	.clk(!CLK),
	.d(\reg_file[30][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][3] .is_wysiwyg = "true";
defparam \reg_file[30][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N9
dffeas \reg_file[18][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][3] .is_wysiwyg = "true";
defparam \reg_file[18][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N10
cycloneive_lcell_comb \reg_file[22][3]~feeder (
// Equation(s):
// \reg_file[22][3]~feeder_combout  = \reg_file_nxt[31][3]~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][3]~66_combout ),
	.cin(gnd),
	.combout(\reg_file[22][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][3]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[22][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N11
dffeas \reg_file[22][3] (
	.clk(!CLK),
	.d(\reg_file[22][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][3] .is_wysiwyg = "true";
defparam \reg_file[22][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N8
cycloneive_lcell_comb \Mux60~2 (
// Equation(s):
// \Mux60~2_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[22][3]~q ))) # (!\prif.imemload_id [18] & (\reg_file[18][3]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][3]~q ),
	.datad(\reg_file[22][3]~q ),
	.cin(gnd),
	.combout(\Mux60~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~2 .lut_mask = 16'hDC98;
defparam \Mux60~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N10
cycloneive_lcell_comb \Mux60~3 (
// Equation(s):
// \Mux60~3_combout  = (\Mux60~2_combout  & (((\reg_file[30][3]~q ) # (!\prif.imemload_id [19])))) # (!\Mux60~2_combout  & (\reg_file[26][3]~q  & ((\prif.imemload_id [19]))))

	.dataa(\reg_file[26][3]~q ),
	.datab(\reg_file[30][3]~q ),
	.datac(\Mux60~2_combout ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux60~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~3 .lut_mask = 16'hCAF0;
defparam \Mux60~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N2
cycloneive_lcell_comb \reg_file[28][3]~feeder (
// Equation(s):
// \reg_file[28][3]~feeder_combout  = \reg_file_nxt[31][3]~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][3]~66_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[28][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[28][3]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[28][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N3
dffeas \reg_file[28][3] (
	.clk(!CLK),
	.d(\reg_file[28][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][3] .is_wysiwyg = "true";
defparam \reg_file[28][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N3
dffeas \reg_file[16][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][3] .is_wysiwyg = "true";
defparam \reg_file[16][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N2
cycloneive_lcell_comb \reg_file[20][3]~feeder (
// Equation(s):
// \reg_file[20][3]~feeder_combout  = \reg_file_nxt[31][3]~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][3]~66_combout ),
	.cin(gnd),
	.combout(\reg_file[20][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[20][3]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[20][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N3
dffeas \reg_file[20][3] (
	.clk(!CLK),
	.d(\reg_file[20][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][3] .is_wysiwyg = "true";
defparam \reg_file[20][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N2
cycloneive_lcell_comb \Mux60~4 (
// Equation(s):
// \Mux60~4_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[20][3]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & (\reg_file[16][3]~q )))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[16][3]~q ),
	.datad(\reg_file[20][3]~q ),
	.cin(gnd),
	.combout(\Mux60~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~4 .lut_mask = 16'hBA98;
defparam \Mux60~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N24
cycloneive_lcell_comb \Mux60~5 (
// Equation(s):
// \Mux60~5_combout  = (\prif.imemload_id [19] & ((\Mux60~4_combout  & ((\reg_file[28][3]~q ))) # (!\Mux60~4_combout  & (\reg_file[24][3]~q )))) # (!\prif.imemload_id [19] & (((\Mux60~4_combout ))))

	.dataa(\reg_file[24][3]~q ),
	.datab(\reg_file[28][3]~q ),
	.datac(prifimemload_id_19),
	.datad(\Mux60~4_combout ),
	.cin(gnd),
	.combout(\Mux60~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~5 .lut_mask = 16'hCFA0;
defparam \Mux60~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N20
cycloneive_lcell_comb \Mux60~6 (
// Equation(s):
// \Mux60~6_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\Mux60~3_combout )) # (!\prif.imemload_id [17] & ((\Mux60~5_combout )))))

	.dataa(\Mux60~3_combout ),
	.datab(prifimemload_id_16),
	.datac(prifimemload_id_17),
	.datad(\Mux60~5_combout ),
	.cin(gnd),
	.combout(\Mux60~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~6 .lut_mask = 16'hE3E0;
defparam \Mux60~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N3
dffeas \reg_file[14][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][3] .is_wysiwyg = "true";
defparam \reg_file[14][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N17
dffeas \reg_file[13][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][3] .is_wysiwyg = "true";
defparam \reg_file[13][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N19
dffeas \reg_file[12][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][3] .is_wysiwyg = "true";
defparam \reg_file[12][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N16
cycloneive_lcell_comb \Mux60~17 (
// Equation(s):
// \Mux60~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & (\reg_file[13][3]~q )) # (!\prif.imemload_id [16] & ((\reg_file[12][3]~q )))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[13][3]~q ),
	.datad(\reg_file[12][3]~q ),
	.cin(gnd),
	.combout(\Mux60~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~17 .lut_mask = 16'hD9C8;
defparam \Mux60~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N29
dffeas \reg_file[15][3] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][3]~66_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][3] .is_wysiwyg = "true";
defparam \reg_file[15][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N10
cycloneive_lcell_comb \Mux60~18 (
// Equation(s):
// \Mux60~18_combout  = (\prif.imemload_id [17] & ((\Mux60~17_combout  & ((\reg_file[15][3]~q ))) # (!\Mux60~17_combout  & (\reg_file[14][3]~q )))) # (!\prif.imemload_id [17] & (((\Mux60~17_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[14][3]~q ),
	.datac(\Mux60~17_combout ),
	.datad(\reg_file[15][3]~q ),
	.cin(gnd),
	.combout(\Mux60~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~18 .lut_mask = 16'hF858;
defparam \Mux60~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y26_N27
dffeas \reg_file[2][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][3] .is_wysiwyg = "true";
defparam \reg_file[2][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N27
dffeas \reg_file[1][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][3] .is_wysiwyg = "true";
defparam \reg_file[1][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N13
dffeas \reg_file[3][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][3] .is_wysiwyg = "true";
defparam \reg_file[3][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N26
cycloneive_lcell_comb \Mux60~14 (
// Equation(s):
// \Mux60~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][3]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][3]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[1][3]~q ),
	.datad(\reg_file[3][3]~q ),
	.cin(gnd),
	.combout(\Mux60~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~14 .lut_mask = 16'hA820;
defparam \Mux60~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N8
cycloneive_lcell_comb \Mux60~15 (
// Equation(s):
// \Mux60~15_combout  = (\Mux60~14_combout ) # ((!\prif.imemload_id [16] & (\reg_file[2][3]~q  & \prif.imemload_id [17])))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[2][3]~q ),
	.datac(\Mux60~14_combout ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux60~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~15 .lut_mask = 16'hF4F0;
defparam \Mux60~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y25_N5
dffeas \reg_file[9][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][3] .is_wysiwyg = "true";
defparam \reg_file[9][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y25_N3
dffeas \reg_file[11][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][3] .is_wysiwyg = "true";
defparam \reg_file[11][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N19
dffeas \reg_file[8][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][3] .is_wysiwyg = "true";
defparam \reg_file[8][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N17
dffeas \reg_file[10][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][3] .is_wysiwyg = "true";
defparam \reg_file[10][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N18
cycloneive_lcell_comb \Mux60~12 (
// Equation(s):
// \Mux60~12_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][3]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][3]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[8][3]~q ),
	.datad(\reg_file[10][3]~q ),
	.cin(gnd),
	.combout(\Mux60~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~12 .lut_mask = 16'hDC98;
defparam \Mux60~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N2
cycloneive_lcell_comb \Mux60~13 (
// Equation(s):
// \Mux60~13_combout  = (\prif.imemload_id [16] & ((\Mux60~12_combout  & ((\reg_file[11][3]~q ))) # (!\Mux60~12_combout  & (\reg_file[9][3]~q )))) # (!\prif.imemload_id [16] & (((\Mux60~12_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[9][3]~q ),
	.datac(\reg_file[11][3]~q ),
	.datad(\Mux60~12_combout ),
	.cin(gnd),
	.combout(\Mux60~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~13 .lut_mask = 16'hF588;
defparam \Mux60~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N30
cycloneive_lcell_comb \Mux60~16 (
// Equation(s):
// \Mux60~16_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18]) # (\Mux60~13_combout )))) # (!\prif.imemload_id [19] & (\Mux60~15_combout  & (!\prif.imemload_id [18])))

	.dataa(prifimemload_id_19),
	.datab(\Mux60~15_combout ),
	.datac(prifimemload_id_18),
	.datad(\Mux60~13_combout ),
	.cin(gnd),
	.combout(\Mux60~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~16 .lut_mask = 16'hAEA4;
defparam \Mux60~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N4
cycloneive_lcell_comb \reg_file[6][3]~feeder (
// Equation(s):
// \reg_file[6][3]~feeder_combout  = \reg_file_nxt[31][3]~66_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][3]~66_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][3]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][3]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][3]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N5
dffeas \reg_file[6][3] (
	.clk(!CLK),
	.d(\reg_file[6][3]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][3] .is_wysiwyg = "true";
defparam \reg_file[6][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y26_N3
dffeas \reg_file[7][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][3] .is_wysiwyg = "true";
defparam \reg_file[7][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N29
dffeas \reg_file[5][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][3] .is_wysiwyg = "true";
defparam \reg_file[5][3] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N11
dffeas \reg_file[4][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][3] .is_wysiwyg = "true";
defparam \reg_file[4][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N28
cycloneive_lcell_comb \Mux60~10 (
// Equation(s):
// \Mux60~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][3]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][3]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][3]~q ),
	.datad(\reg_file[4][3]~q ),
	.cin(gnd),
	.combout(\Mux60~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~10 .lut_mask = 16'hB9A8;
defparam \Mux60~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N16
cycloneive_lcell_comb \Mux60~11 (
// Equation(s):
// \Mux60~11_combout  = (\prif.imemload_id [17] & ((\Mux60~10_combout  & ((\reg_file[7][3]~q ))) # (!\Mux60~10_combout  & (\reg_file[6][3]~q )))) # (!\prif.imemload_id [17] & (((\Mux60~10_combout ))))

	.dataa(\reg_file[6][3]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[7][3]~q ),
	.datad(\Mux60~10_combout ),
	.cin(gnd),
	.combout(\Mux60~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux60~11 .lut_mask = 16'hF388;
defparam \Mux60~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N22
cycloneive_lcell_comb \reg_file_nxt[31][2]~67 (
// Equation(s):
// \reg_file_nxt[31][2]~67_combout  = (\Mux162~1_combout  & ((\prif.regwrite_wb [0]) # ((\prif.regwrite_wb [2]) # (!Equal8))))

	.dataa(Mux162),
	.datab(prifregwrite_wb_0),
	.datac(Equal8),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\reg_file_nxt[31][2]~67_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][2]~67 .lut_mask = 16'hAA8A;
defparam \reg_file_nxt[31][2]~67 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N21
dffeas \reg_file[22][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][2] .is_wysiwyg = "true";
defparam \reg_file[22][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N24
cycloneive_lcell_comb \reg_file[18][2]~feeder (
// Equation(s):
// \reg_file[18][2]~feeder_combout  = \reg_file_nxt[31][2]~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][2]~67_combout ),
	.cin(gnd),
	.combout(\reg_file[18][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[18][2]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[18][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y30_N25
dffeas \reg_file[18][2] (
	.clk(!CLK),
	.d(\reg_file[18][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][2] .is_wysiwyg = "true";
defparam \reg_file[18][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N24
cycloneive_lcell_comb \reg_file[26][2]~feeder (
// Equation(s):
// \reg_file[26][2]~feeder_combout  = \reg_file_nxt[31][2]~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][2]~67_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[26][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[26][2]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[26][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N25
dffeas \reg_file[26][2] (
	.clk(!CLK),
	.d(\reg_file[26][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][2] .is_wysiwyg = "true";
defparam \reg_file[26][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N30
cycloneive_lcell_comb \Mux61~2 (
// Equation(s):
// \Mux61~2_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18]) # (\reg_file[26][2]~q )))) # (!\prif.imemload_id [19] & (\reg_file[18][2]~q  & (!\prif.imemload_id [18])))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[18][2]~q ),
	.datac(prifimemload_id_18),
	.datad(\reg_file[26][2]~q ),
	.cin(gnd),
	.combout(\Mux61~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~2 .lut_mask = 16'hAEA4;
defparam \Mux61~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N28
cycloneive_lcell_comb \Mux61~3 (
// Equation(s):
// \Mux61~3_combout  = (\prif.imemload_id [18] & ((\Mux61~2_combout  & (\reg_file[30][2]~q )) # (!\Mux61~2_combout  & ((\reg_file[22][2]~q ))))) # (!\prif.imemload_id [18] & (((\Mux61~2_combout ))))

	.dataa(\reg_file[30][2]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[22][2]~q ),
	.datad(\Mux61~2_combout ),
	.cin(gnd),
	.combout(\Mux61~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~3 .lut_mask = 16'hBBC0;
defparam \Mux61~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N21
dffeas \reg_file[20][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][2] .is_wysiwyg = "true";
defparam \reg_file[20][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y33_N1
dffeas \reg_file[24][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][2] .is_wysiwyg = "true";
defparam \reg_file[24][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N0
cycloneive_lcell_comb \Mux61~4 (
// Equation(s):
// \Mux61~4_combout  = (\prif.imemload_id [19] & (((\reg_file[24][2]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[16][2]~q  & ((!\prif.imemload_id [18]))))

	.dataa(\reg_file[16][2]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[24][2]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux61~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~4 .lut_mask = 16'hCCE2;
defparam \Mux61~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N20
cycloneive_lcell_comb \Mux61~5 (
// Equation(s):
// \Mux61~5_combout  = (\prif.imemload_id [18] & ((\Mux61~4_combout  & (\reg_file[28][2]~q )) # (!\Mux61~4_combout  & ((\reg_file[20][2]~q ))))) # (!\prif.imemload_id [18] & (((\Mux61~4_combout ))))

	.dataa(\reg_file[28][2]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[20][2]~q ),
	.datad(\Mux61~4_combout ),
	.cin(gnd),
	.combout(\Mux61~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~5 .lut_mask = 16'hBBC0;
defparam \Mux61~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N6
cycloneive_lcell_comb \Mux61~6 (
// Equation(s):
// \Mux61~6_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\Mux61~3_combout )) # (!\prif.imemload_id [17] & ((\Mux61~5_combout )))))

	.dataa(prifimemload_id_16),
	.datab(\Mux61~3_combout ),
	.datac(prifimemload_id_17),
	.datad(\Mux61~5_combout ),
	.cin(gnd),
	.combout(\Mux61~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~6 .lut_mask = 16'hE5E0;
defparam \Mux61~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N29
dffeas \reg_file[23][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][2] .is_wysiwyg = "true";
defparam \reg_file[23][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N21
dffeas \reg_file[19][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][2] .is_wysiwyg = "true";
defparam \reg_file[19][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N28
cycloneive_lcell_comb \Mux61~7 (
// Equation(s):
// \Mux61~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][2]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][2]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][2]~q ),
	.datad(\reg_file[19][2]~q ),
	.cin(gnd),
	.combout(\Mux61~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~7 .lut_mask = 16'hB9A8;
defparam \Mux61~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N22
cycloneive_lcell_comb \reg_file[31][2]~feeder (
// Equation(s):
// \reg_file[31][2]~feeder_combout  = \reg_file_nxt[31][2]~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][2]~67_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[31][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][2]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[31][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y27_N23
dffeas \reg_file[31][2] (
	.clk(!CLK),
	.d(\reg_file[31][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][2] .is_wysiwyg = "true";
defparam \reg_file[31][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N22
cycloneive_lcell_comb \reg_file[27][2]~feeder (
// Equation(s):
// \reg_file[27][2]~feeder_combout  = \reg_file_nxt[31][2]~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][2]~67_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[27][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[27][2]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[27][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N23
dffeas \reg_file[27][2] (
	.clk(!CLK),
	.d(\reg_file[27][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][2] .is_wysiwyg = "true";
defparam \reg_file[27][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N28
cycloneive_lcell_comb \Mux61~8 (
// Equation(s):
// \Mux61~8_combout  = (\prif.imemload_id [19] & ((\Mux61~7_combout  & (\reg_file[31][2]~q )) # (!\Mux61~7_combout  & ((\reg_file[27][2]~q ))))) # (!\prif.imemload_id [19] & (\Mux61~7_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux61~7_combout ),
	.datac(\reg_file[31][2]~q ),
	.datad(\reg_file[27][2]~q ),
	.cin(gnd),
	.combout(\Mux61~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~8 .lut_mask = 16'hE6C4;
defparam \Mux61~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N3
dffeas \reg_file[25][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][2] .is_wysiwyg = "true";
defparam \reg_file[25][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N2
cycloneive_lcell_comb \reg_file[29][2]~feeder (
// Equation(s):
// \reg_file[29][2]~feeder_combout  = \reg_file_nxt[31][2]~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][2]~67_combout ),
	.cin(gnd),
	.combout(\reg_file[29][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][2]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N3
dffeas \reg_file[29][2] (
	.clk(!CLK),
	.d(\reg_file[29][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][2] .is_wysiwyg = "true";
defparam \reg_file[29][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N17
dffeas \reg_file[17][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][2] .is_wysiwyg = "true";
defparam \reg_file[17][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y24_N16
cycloneive_lcell_comb \reg_file[21][2]~feeder (
// Equation(s):
// \reg_file[21][2]~feeder_combout  = \reg_file_nxt[31][2]~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][2]~67_combout ),
	.cin(gnd),
	.combout(\reg_file[21][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][2]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[21][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y24_N17
dffeas \reg_file[21][2] (
	.clk(!CLK),
	.d(\reg_file[21][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][2] .is_wysiwyg = "true";
defparam \reg_file[21][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N16
cycloneive_lcell_comb \Mux61~0 (
// Equation(s):
// \Mux61~0_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[21][2]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & (\reg_file[17][2]~q )))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][2]~q ),
	.datad(\reg_file[21][2]~q ),
	.cin(gnd),
	.combout(\Mux61~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~0 .lut_mask = 16'hBA98;
defparam \Mux61~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N28
cycloneive_lcell_comb \Mux61~1 (
// Equation(s):
// \Mux61~1_combout  = (\prif.imemload_id [19] & ((\Mux61~0_combout  & ((\reg_file[29][2]~q ))) # (!\Mux61~0_combout  & (\reg_file[25][2]~q )))) # (!\prif.imemload_id [19] & (((\Mux61~0_combout ))))

	.dataa(\reg_file[25][2]~q ),
	.datab(\reg_file[29][2]~q ),
	.datac(prifimemload_id_19),
	.datad(\Mux61~0_combout ),
	.cin(gnd),
	.combout(\Mux61~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~1 .lut_mask = 16'hCFA0;
defparam \Mux61~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y25_N9
dffeas \reg_file[10][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][2] .is_wysiwyg = "true";
defparam \reg_file[10][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N8
cycloneive_lcell_comb \Mux61~10 (
// Equation(s):
// \Mux61~10_combout  = (\prif.imemload_id [17] & (((\reg_file[10][2]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][2]~q  & ((!\prif.imemload_id [16]))))

	.dataa(\reg_file[8][2]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[10][2]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux61~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~10 .lut_mask = 16'hCCE2;
defparam \Mux61~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y25_N29
dffeas \reg_file[9][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][2] .is_wysiwyg = "true";
defparam \reg_file[9][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y25_N11
dffeas \reg_file[11][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][2] .is_wysiwyg = "true";
defparam \reg_file[11][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N28
cycloneive_lcell_comb \Mux61~11 (
// Equation(s):
// \Mux61~11_combout  = (\prif.imemload_id [16] & ((\Mux61~10_combout  & ((\reg_file[11][2]~q ))) # (!\Mux61~10_combout  & (\reg_file[9][2]~q )))) # (!\prif.imemload_id [16] & (\Mux61~10_combout ))

	.dataa(prifimemload_id_16),
	.datab(\Mux61~10_combout ),
	.datac(\reg_file[9][2]~q ),
	.datad(\reg_file[11][2]~q ),
	.cin(gnd),
	.combout(\Mux61~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~11 .lut_mask = 16'hEC64;
defparam \Mux61~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N23
dffeas \reg_file[15][2] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][2]~67_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][2] .is_wysiwyg = "true";
defparam \reg_file[15][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y26_N13
dffeas \reg_file[14][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][2] .is_wysiwyg = "true";
defparam \reg_file[14][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N15
dffeas \reg_file[12][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][2] .is_wysiwyg = "true";
defparam \reg_file[12][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N25
dffeas \reg_file[13][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][2] .is_wysiwyg = "true";
defparam \reg_file[13][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N14
cycloneive_lcell_comb \Mux61~17 (
// Equation(s):
// \Mux61~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][2]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][2]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][2]~q ),
	.datad(\reg_file[13][2]~q ),
	.cin(gnd),
	.combout(\Mux61~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~17 .lut_mask = 16'hDC98;
defparam \Mux61~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N8
cycloneive_lcell_comb \Mux61~18 (
// Equation(s):
// \Mux61~18_combout  = (\prif.imemload_id [17] & ((\Mux61~17_combout  & (\reg_file[15][2]~q )) # (!\Mux61~17_combout  & ((\reg_file[14][2]~q ))))) # (!\prif.imemload_id [17] & (((\Mux61~17_combout ))))

	.dataa(\reg_file[15][2]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[14][2]~q ),
	.datad(\Mux61~17_combout ),
	.cin(gnd),
	.combout(\Mux61~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~18 .lut_mask = 16'hBBC0;
defparam \Mux61~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y27_N3
dffeas \reg_file[7][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][2] .is_wysiwyg = "true";
defparam \reg_file[7][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N11
dffeas \reg_file[4][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][2] .is_wysiwyg = "true";
defparam \reg_file[4][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N13
dffeas \reg_file[5][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][2] .is_wysiwyg = "true";
defparam \reg_file[5][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N10
cycloneive_lcell_comb \Mux61~12 (
// Equation(s):
// \Mux61~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][2]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][2]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][2]~q ),
	.datad(\reg_file[5][2]~q ),
	.cin(gnd),
	.combout(\Mux61~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~12 .lut_mask = 16'hBA98;
defparam \Mux61~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N2
cycloneive_lcell_comb \Mux61~13 (
// Equation(s):
// \Mux61~13_combout  = (\prif.imemload_id [17] & ((\Mux61~12_combout  & ((\reg_file[7][2]~q ))) # (!\Mux61~12_combout  & (\reg_file[6][2]~q )))) # (!\prif.imemload_id [17] & (((\Mux61~12_combout ))))

	.dataa(\reg_file[6][2]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[7][2]~q ),
	.datad(\Mux61~12_combout ),
	.cin(gnd),
	.combout(\Mux61~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~13 .lut_mask = 16'hF388;
defparam \Mux61~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y27_N1
dffeas \reg_file[2][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][2] .is_wysiwyg = "true";
defparam \reg_file[2][2] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y25_N15
dffeas \reg_file[1][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][2] .is_wysiwyg = "true";
defparam \reg_file[1][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N12
cycloneive_lcell_comb \reg_file[3][2]~feeder (
// Equation(s):
// \reg_file[3][2]~feeder_combout  = \reg_file_nxt[31][2]~67_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][2]~67_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[3][2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[3][2]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[3][2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y25_N13
dffeas \reg_file[3][2] (
	.clk(!CLK),
	.d(\reg_file[3][2]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][2] .is_wysiwyg = "true";
defparam \reg_file[3][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N14
cycloneive_lcell_comb \Mux61~14 (
// Equation(s):
// \Mux61~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][2]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][2]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[1][2]~q ),
	.datad(\reg_file[3][2]~q ),
	.cin(gnd),
	.combout(\Mux61~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~14 .lut_mask = 16'hA820;
defparam \Mux61~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N0
cycloneive_lcell_comb \Mux61~15 (
// Equation(s):
// \Mux61~15_combout  = (\Mux61~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][2]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[2][2]~q ),
	.datad(\Mux61~14_combout ),
	.cin(gnd),
	.combout(\Mux61~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~15 .lut_mask = 16'hFF40;
defparam \Mux61~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N10
cycloneive_lcell_comb \Mux61~16 (
// Equation(s):
// \Mux61~16_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\Mux61~13_combout )) # (!\prif.imemload_id [18] & ((\Mux61~15_combout )))))

	.dataa(prifimemload_id_19),
	.datab(\Mux61~13_combout ),
	.datac(prifimemload_id_18),
	.datad(\Mux61~15_combout ),
	.cin(gnd),
	.combout(\Mux61~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux61~16 .lut_mask = 16'hE5E0;
defparam \Mux61~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N26
cycloneive_lcell_comb \reg_file_nxt[31][4]~68 (
// Equation(s):
// \reg_file_nxt[31][4]~68_combout  = (\Mux160~1_combout  & ((\prif.regwrite_wb [0]) # ((\prif.regwrite_wb [2]) # (!Equal8))))

	.dataa(Mux160),
	.datab(prifregwrite_wb_0),
	.datac(Equal8),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\reg_file_nxt[31][4]~68_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][4]~68 .lut_mask = 16'hAA8A;
defparam \reg_file_nxt[31][4]~68 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N30
cycloneive_lcell_comb \reg_file[27][4]~feeder (
// Equation(s):
// \reg_file[27][4]~feeder_combout  = \reg_file_nxt[31][4]~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][4]~68_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[27][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[27][4]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[27][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N31
dffeas \reg_file[27][4] (
	.clk(!CLK),
	.d(\reg_file[27][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][4] .is_wysiwyg = "true";
defparam \reg_file[27][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N21
dffeas \reg_file[23][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][4] .is_wysiwyg = "true";
defparam \reg_file[23][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N31
dffeas \reg_file[19][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][4] .is_wysiwyg = "true";
defparam \reg_file[19][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N20
cycloneive_lcell_comb \Mux59~7 (
// Equation(s):
// \Mux59~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][4]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][4]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][4]~q ),
	.datad(\reg_file[19][4]~q ),
	.cin(gnd),
	.combout(\Mux59~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~7 .lut_mask = 16'hB9A8;
defparam \Mux59~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y27_N5
dffeas \reg_file[31][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][4] .is_wysiwyg = "true";
defparam \reg_file[31][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N4
cycloneive_lcell_comb \Mux59~8 (
// Equation(s):
// \Mux59~8_combout  = (\Mux59~7_combout  & (((\reg_file[31][4]~q ) # (!\prif.imemload_id [19])))) # (!\Mux59~7_combout  & (\reg_file[27][4]~q  & ((\prif.imemload_id [19]))))

	.dataa(\reg_file[27][4]~q ),
	.datab(\Mux59~7_combout ),
	.datac(\reg_file[31][4]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux59~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~8 .lut_mask = 16'hE2CC;
defparam \Mux59~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N4
cycloneive_lcell_comb \reg_file[22][4]~feeder (
// Equation(s):
// \reg_file[22][4]~feeder_combout  = \reg_file_nxt[31][4]~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][4]~68_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[22][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][4]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[22][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N5
dffeas \reg_file[22][4] (
	.clk(!CLK),
	.d(\reg_file[22][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][4] .is_wysiwyg = "true";
defparam \reg_file[22][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N3
dffeas \reg_file[30][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][4] .is_wysiwyg = "true";
defparam \reg_file[30][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N29
dffeas \reg_file[26][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][4] .is_wysiwyg = "true";
defparam \reg_file[26][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N5
dffeas \reg_file[18][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][4] .is_wysiwyg = "true";
defparam \reg_file[18][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N4
cycloneive_lcell_comb \Mux59~2 (
// Equation(s):
// \Mux59~2_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[26][4]~q )) # (!\prif.imemload_id [19] & ((\reg_file[18][4]~q )))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[26][4]~q ),
	.datac(\reg_file[18][4]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux59~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~2 .lut_mask = 16'hEE50;
defparam \Mux59~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N2
cycloneive_lcell_comb \Mux59~3 (
// Equation(s):
// \Mux59~3_combout  = (\prif.imemload_id [18] & ((\Mux59~2_combout  & ((\reg_file[30][4]~q ))) # (!\Mux59~2_combout  & (\reg_file[22][4]~q )))) # (!\prif.imemload_id [18] & (((\Mux59~2_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[22][4]~q ),
	.datac(\reg_file[30][4]~q ),
	.datad(\Mux59~2_combout ),
	.cin(gnd),
	.combout(\Mux59~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~3 .lut_mask = 16'hF588;
defparam \Mux59~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N7
dffeas \reg_file[28][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][4] .is_wysiwyg = "true";
defparam \reg_file[28][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N25
dffeas \reg_file[20][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][4] .is_wysiwyg = "true";
defparam \reg_file[20][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N24
cycloneive_lcell_comb \Mux59~5 (
// Equation(s):
// \Mux59~5_combout  = (\Mux59~4_combout  & ((\reg_file[28][4]~q ) # ((!\prif.imemload_id [18])))) # (!\Mux59~4_combout  & (((\reg_file[20][4]~q  & \prif.imemload_id [18]))))

	.dataa(\Mux59~4_combout ),
	.datab(\reg_file[28][4]~q ),
	.datac(\reg_file[20][4]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux59~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~5 .lut_mask = 16'hD8AA;
defparam \Mux59~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y27_N4
cycloneive_lcell_comb \Mux59~6 (
// Equation(s):
// \Mux59~6_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\Mux59~3_combout )) # (!\prif.imemload_id [17] & ((\Mux59~5_combout )))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\Mux59~3_combout ),
	.datad(\Mux59~5_combout ),
	.cin(gnd),
	.combout(\Mux59~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~6 .lut_mask = 16'hD9C8;
defparam \Mux59~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N12
cycloneive_lcell_comb \reg_file[29][4]~feeder (
// Equation(s):
// \reg_file[29][4]~feeder_combout  = \reg_file_nxt[31][4]~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][4]~68_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][4]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N13
dffeas \reg_file[29][4] (
	.clk(!CLK),
	.d(\reg_file[29][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][4] .is_wysiwyg = "true";
defparam \reg_file[29][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N23
dffeas \reg_file[17][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][4] .is_wysiwyg = "true";
defparam \reg_file[17][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y24_N2
cycloneive_lcell_comb \reg_file[21][4]~feeder (
// Equation(s):
// \reg_file[21][4]~feeder_combout  = \reg_file_nxt[31][4]~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][4]~68_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[21][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][4]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[21][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y24_N3
dffeas \reg_file[21][4] (
	.clk(!CLK),
	.d(\reg_file[21][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][4] .is_wysiwyg = "true";
defparam \reg_file[21][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N22
cycloneive_lcell_comb \Mux59~0 (
// Equation(s):
// \Mux59~0_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[21][4]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & (\reg_file[17][4]~q )))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][4]~q ),
	.datad(\reg_file[21][4]~q ),
	.cin(gnd),
	.combout(\Mux59~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~0 .lut_mask = 16'hBA98;
defparam \Mux59~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N31
dffeas \reg_file[25][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][4] .is_wysiwyg = "true";
defparam \reg_file[25][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N22
cycloneive_lcell_comb \Mux59~1 (
// Equation(s):
// \Mux59~1_combout  = (\Mux59~0_combout  & ((\reg_file[29][4]~q ) # ((!\prif.imemload_id [19])))) # (!\Mux59~0_combout  & (((\reg_file[25][4]~q  & \prif.imemload_id [19]))))

	.dataa(\reg_file[29][4]~q ),
	.datab(\Mux59~0_combout ),
	.datac(\reg_file[25][4]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux59~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~1 .lut_mask = 16'hB8CC;
defparam \Mux59~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y25_N21
dffeas \reg_file[10][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][4] .is_wysiwyg = "true";
defparam \reg_file[10][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N20
cycloneive_lcell_comb \Mux59~10 (
// Equation(s):
// \Mux59~10_combout  = (\prif.imemload_id [17] & (((\reg_file[10][4]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][4]~q  & ((!\prif.imemload_id [16]))))

	.dataa(\reg_file[8][4]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[10][4]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux59~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~10 .lut_mask = 16'hCCE2;
defparam \Mux59~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y25_N17
dffeas \reg_file[9][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][4] .is_wysiwyg = "true";
defparam \reg_file[9][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y25_N7
dffeas \reg_file[11][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][4] .is_wysiwyg = "true";
defparam \reg_file[11][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N16
cycloneive_lcell_comb \Mux59~11 (
// Equation(s):
// \Mux59~11_combout  = (\prif.imemload_id [16] & ((\Mux59~10_combout  & ((\reg_file[11][4]~q ))) # (!\Mux59~10_combout  & (\reg_file[9][4]~q )))) # (!\prif.imemload_id [16] & (\Mux59~10_combout ))

	.dataa(prifimemload_id_16),
	.datab(\Mux59~10_combout ),
	.datac(\reg_file[9][4]~q ),
	.datad(\reg_file[11][4]~q ),
	.cin(gnd),
	.combout(\Mux59~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~11 .lut_mask = 16'hEC64;
defparam \Mux59~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y26_N31
dffeas \reg_file[4][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][4] .is_wysiwyg = "true";
defparam \reg_file[4][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N25
dffeas \reg_file[5][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][4] .is_wysiwyg = "true";
defparam \reg_file[5][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N30
cycloneive_lcell_comb \Mux59~12 (
// Equation(s):
// \Mux59~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][4]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][4]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][4]~q ),
	.datad(\reg_file[5][4]~q ),
	.cin(gnd),
	.combout(\Mux59~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~12 .lut_mask = 16'hBA98;
defparam \Mux59~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y25_N25
dffeas \reg_file[7][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][4] .is_wysiwyg = "true";
defparam \reg_file[7][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N30
cycloneive_lcell_comb \Mux59~13 (
// Equation(s):
// \Mux59~13_combout  = (\Mux59~12_combout  & (((\reg_file[7][4]~q ) # (!\prif.imemload_id [17])))) # (!\Mux59~12_combout  & (\reg_file[6][4]~q  & (\prif.imemload_id [17])))

	.dataa(\reg_file[6][4]~q ),
	.datab(\Mux59~12_combout ),
	.datac(prifimemload_id_17),
	.datad(\reg_file[7][4]~q ),
	.cin(gnd),
	.combout(\Mux59~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~13 .lut_mask = 16'hEC2C;
defparam \Mux59~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N20
cycloneive_lcell_comb \reg_file[2][4]~feeder (
// Equation(s):
// \reg_file[2][4]~feeder_combout  = \reg_file_nxt[31][4]~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][4]~68_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[2][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][4]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[2][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y25_N21
dffeas \reg_file[2][4] (
	.clk(!CLK),
	.d(\reg_file[2][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][4] .is_wysiwyg = "true";
defparam \reg_file[2][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y25_N29
dffeas \reg_file[1][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][4] .is_wysiwyg = "true";
defparam \reg_file[1][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N28
cycloneive_lcell_comb \Mux59~14 (
// Equation(s):
// \Mux59~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][4]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][4]~q )))))

	.dataa(\reg_file[3][4]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[1][4]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux59~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~14 .lut_mask = 16'hB800;
defparam \Mux59~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N6
cycloneive_lcell_comb \Mux59~15 (
// Equation(s):
// \Mux59~15_combout  = (\Mux59~14_combout ) # ((!\prif.imemload_id [16] & (\reg_file[2][4]~q  & \prif.imemload_id [17])))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[2][4]~q ),
	.datac(prifimemload_id_17),
	.datad(\Mux59~14_combout ),
	.cin(gnd),
	.combout(\Mux59~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~15 .lut_mask = 16'hFF40;
defparam \Mux59~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N4
cycloneive_lcell_comb \Mux59~16 (
// Equation(s):
// \Mux59~16_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\Mux59~13_combout )) # (!\prif.imemload_id [18] & ((\Mux59~15_combout )))))

	.dataa(\Mux59~13_combout ),
	.datab(prifimemload_id_19),
	.datac(prifimemload_id_18),
	.datad(\Mux59~15_combout ),
	.cin(gnd),
	.combout(\Mux59~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~16 .lut_mask = 16'hE3E0;
defparam \Mux59~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N21
dffeas \reg_file[14][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][4] .is_wysiwyg = "true";
defparam \reg_file[14][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N23
dffeas \reg_file[12][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][4] .is_wysiwyg = "true";
defparam \reg_file[12][4] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N21
dffeas \reg_file[13][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][4] .is_wysiwyg = "true";
defparam \reg_file[13][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N22
cycloneive_lcell_comb \Mux59~17 (
// Equation(s):
// \Mux59~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][4]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][4]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][4]~q ),
	.datad(\reg_file[13][4]~q ),
	.cin(gnd),
	.combout(\Mux59~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~17 .lut_mask = 16'hDC98;
defparam \Mux59~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N27
dffeas \reg_file[15][4] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][4]~68_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][4] .is_wysiwyg = "true";
defparam \reg_file[15][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N2
cycloneive_lcell_comb \Mux59~18 (
// Equation(s):
// \Mux59~18_combout  = (\Mux59~17_combout  & (((\reg_file[15][4]~q ) # (!\prif.imemload_id [17])))) # (!\Mux59~17_combout  & (\reg_file[14][4]~q  & ((\prif.imemload_id [17]))))

	.dataa(\reg_file[14][4]~q ),
	.datab(\Mux59~17_combout ),
	.datac(\reg_file[15][4]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux59~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux59~18 .lut_mask = 16'hE2CC;
defparam \Mux59~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N14
cycloneive_lcell_comb \reg_file_nxt[31][31]~69 (
// Equation(s):
// \reg_file_nxt[31][31]~69_combout  = (\Mux133~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(Mux133),
	.datab(prifregwrite_wb_2),
	.datac(Equal8),
	.datad(prifregwrite_wb_0),
	.cin(gnd),
	.combout(\reg_file_nxt[31][31]~69_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][31]~69 .lut_mask = 16'hAA8A;
defparam \reg_file_nxt[31][31]~69 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N21
dffeas \reg_file[21][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][31] .is_wysiwyg = "true";
defparam \reg_file[21][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N14
cycloneive_lcell_comb \reg_file[29][31]~feeder (
// Equation(s):
// \reg_file[29][31]~feeder_combout  = \reg_file_nxt[31][31]~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][31]~69_combout ),
	.cin(gnd),
	.combout(\reg_file[29][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][31]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N15
dffeas \reg_file[29][31] (
	.clk(!CLK),
	.d(\reg_file[29][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][31] .is_wysiwyg = "true";
defparam \reg_file[29][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N21
dffeas \reg_file[17][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][31] .is_wysiwyg = "true";
defparam \reg_file[17][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N28
cycloneive_lcell_comb \reg_file[25][31]~feeder (
// Equation(s):
// \reg_file[25][31]~feeder_combout  = \reg_file_nxt[31][31]~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][31]~69_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[25][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][31]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[25][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N29
dffeas \reg_file[25][31] (
	.clk(!CLK),
	.d(\reg_file[25][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][31] .is_wysiwyg = "true";
defparam \reg_file[25][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N20
cycloneive_lcell_comb \Mux32~0 (
// Equation(s):
// \Mux32~0_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[25][31]~q ))) # (!\prif.imemload_id [19] & (\reg_file[17][31]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][31]~q ),
	.datad(\reg_file[25][31]~q ),
	.cin(gnd),
	.combout(\Mux32~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~0 .lut_mask = 16'hDC98;
defparam \Mux32~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N28
cycloneive_lcell_comb \Mux32~1 (
// Equation(s):
// \Mux32~1_combout  = (\prif.imemload_id [18] & ((\Mux32~0_combout  & ((\reg_file[29][31]~q ))) # (!\Mux32~0_combout  & (\reg_file[21][31]~q )))) # (!\prif.imemload_id [18] & (((\Mux32~0_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[21][31]~q ),
	.datac(\reg_file[29][31]~q ),
	.datad(\Mux32~0_combout ),
	.cin(gnd),
	.combout(\Mux32~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~1 .lut_mask = 16'hF588;
defparam \Mux32~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N9
dffeas \reg_file[24][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][31] .is_wysiwyg = "true";
defparam \reg_file[24][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N2
cycloneive_lcell_comb \reg_file[28][31]~feeder (
// Equation(s):
// \reg_file[28][31]~feeder_combout  = \reg_file_nxt[31][31]~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][31]~69_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[28][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[28][31]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[28][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N3
dffeas \reg_file[28][31] (
	.clk(!CLK),
	.d(\reg_file[28][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][31] .is_wysiwyg = "true";
defparam \reg_file[28][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N8
cycloneive_lcell_comb \Mux32~5 (
// Equation(s):
// \Mux32~5_combout  = (\Mux32~4_combout  & (((\reg_file[28][31]~q )) # (!\prif.imemload_id [19]))) # (!\Mux32~4_combout  & (\prif.imemload_id [19] & (\reg_file[24][31]~q )))

	.dataa(\Mux32~4_combout ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[24][31]~q ),
	.datad(\reg_file[28][31]~q ),
	.cin(gnd),
	.combout(\Mux32~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~5 .lut_mask = 16'hEA62;
defparam \Mux32~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y30_N19
dffeas \reg_file[18][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][31] .is_wysiwyg = "true";
defparam \reg_file[18][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N18
cycloneive_lcell_comb \Mux32~2 (
// Equation(s):
// \Mux32~2_combout  = (\prif.imemload_id [18] & ((\reg_file[22][31]~q ) # ((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (((\reg_file[18][31]~q  & !\prif.imemload_id [19]))))

	.dataa(\reg_file[22][31]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][31]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux32~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~2 .lut_mask = 16'hCCB8;
defparam \Mux32~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N7
dffeas \reg_file[30][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][31] .is_wysiwyg = "true";
defparam \reg_file[30][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N19
dffeas \reg_file[26][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][31] .is_wysiwyg = "true";
defparam \reg_file[26][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N6
cycloneive_lcell_comb \Mux32~3 (
// Equation(s):
// \Mux32~3_combout  = (\prif.imemload_id [19] & ((\Mux32~2_combout  & (\reg_file[30][31]~q )) # (!\Mux32~2_combout  & ((\reg_file[26][31]~q ))))) # (!\prif.imemload_id [19] & (\Mux32~2_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux32~2_combout ),
	.datac(\reg_file[30][31]~q ),
	.datad(\reg_file[26][31]~q ),
	.cin(gnd),
	.combout(\Mux32~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~3 .lut_mask = 16'hE6C4;
defparam \Mux32~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N26
cycloneive_lcell_comb \Mux32~6 (
// Equation(s):
// \Mux32~6_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16]) # (\Mux32~3_combout )))) # (!\prif.imemload_id [17] & (\Mux32~5_combout  & (!\prif.imemload_id [16])))

	.dataa(prifimemload_id_17),
	.datab(\Mux32~5_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux32~3_combout ),
	.cin(gnd),
	.combout(\Mux32~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~6 .lut_mask = 16'hAEA4;
defparam \Mux32~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N22
cycloneive_lcell_comb \reg_file[23][31]~feeder (
// Equation(s):
// \reg_file[23][31]~feeder_combout  = \reg_file_nxt[31][31]~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][31]~69_combout ),
	.cin(gnd),
	.combout(\reg_file[23][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][31]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[23][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N23
dffeas \reg_file[23][31] (
	.clk(!CLK),
	.d(\reg_file[23][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][31] .is_wysiwyg = "true";
defparam \reg_file[23][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y26_N17
dffeas \reg_file[27][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][31] .is_wysiwyg = "true";
defparam \reg_file[27][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N9
dffeas \reg_file[19][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][31] .is_wysiwyg = "true";
defparam \reg_file[19][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N16
cycloneive_lcell_comb \Mux32~7 (
// Equation(s):
// \Mux32~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][31]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][31]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][31]~q ),
	.datad(\reg_file[19][31]~q ),
	.cin(gnd),
	.combout(\Mux32~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~7 .lut_mask = 16'hD9C8;
defparam \Mux32~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y26_N23
dffeas \reg_file[31][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][31] .is_wysiwyg = "true";
defparam \reg_file[31][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N14
cycloneive_lcell_comb \Mux32~8 (
// Equation(s):
// \Mux32~8_combout  = (\Mux32~7_combout  & (((\reg_file[31][31]~q ) # (!\prif.imemload_id [18])))) # (!\Mux32~7_combout  & (\reg_file[23][31]~q  & ((\prif.imemload_id [18]))))

	.dataa(\reg_file[23][31]~q ),
	.datab(\Mux32~7_combout ),
	.datac(\reg_file[31][31]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux32~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~8 .lut_mask = 16'hE2CC;
defparam \Mux32~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N25
dffeas \reg_file[14][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][31] .is_wysiwyg = "true";
defparam \reg_file[14][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y26_N15
dffeas \reg_file[15][31] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][31]~69_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][31] .is_wysiwyg = "true";
defparam \reg_file[15][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N7
dffeas \reg_file[12][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][31] .is_wysiwyg = "true";
defparam \reg_file[12][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N25
dffeas \reg_file[13][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][31] .is_wysiwyg = "true";
defparam \reg_file[13][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N6
cycloneive_lcell_comb \Mux32~17 (
// Equation(s):
// \Mux32~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][31]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][31]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][31]~q ),
	.datad(\reg_file[13][31]~q ),
	.cin(gnd),
	.combout(\Mux32~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~17 .lut_mask = 16'hDC98;
defparam \Mux32~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N10
cycloneive_lcell_comb \Mux32~18 (
// Equation(s):
// \Mux32~18_combout  = (\prif.imemload_id [17] & ((\Mux32~17_combout  & ((\reg_file[15][31]~q ))) # (!\Mux32~17_combout  & (\reg_file[14][31]~q )))) # (!\prif.imemload_id [17] & (((\Mux32~17_combout ))))

	.dataa(\reg_file[14][31]~q ),
	.datab(\reg_file[15][31]~q ),
	.datac(prifimemload_id_17),
	.datad(\Mux32~17_combout ),
	.cin(gnd),
	.combout(\Mux32~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~18 .lut_mask = 16'hCFA0;
defparam \Mux32~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N15
dffeas \reg_file[7][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][31] .is_wysiwyg = "true";
defparam \reg_file[7][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N23
dffeas \reg_file[4][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][31] .is_wysiwyg = "true";
defparam \reg_file[4][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N23
dffeas \reg_file[5][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][31] .is_wysiwyg = "true";
defparam \reg_file[5][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N22
cycloneive_lcell_comb \Mux32~10 (
// Equation(s):
// \Mux32~10_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[5][31]~q ))) # (!\prif.imemload_id [16] & (\reg_file[4][31]~q ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[4][31]~q ),
	.datac(\reg_file[5][31]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux32~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~10 .lut_mask = 16'hFA44;
defparam \Mux32~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N28
cycloneive_lcell_comb \reg_file[6][31]~feeder (
// Equation(s):
// \reg_file[6][31]~feeder_combout  = \reg_file_nxt[31][31]~69_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][31]~69_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][31]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][31]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][31]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N29
dffeas \reg_file[6][31] (
	.clk(!CLK),
	.d(\reg_file[6][31]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][31] .is_wysiwyg = "true";
defparam \reg_file[6][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y25_N8
cycloneive_lcell_comb \Mux32~11 (
// Equation(s):
// \Mux32~11_combout  = (\prif.imemload_id [17] & ((\Mux32~10_combout  & (\reg_file[7][31]~q )) # (!\Mux32~10_combout  & ((\reg_file[6][31]~q ))))) # (!\prif.imemload_id [17] & (((\Mux32~10_combout ))))

	.dataa(\reg_file[7][31]~q ),
	.datab(prifimemload_id_17),
	.datac(\Mux32~10_combout ),
	.datad(\reg_file[6][31]~q ),
	.cin(gnd),
	.combout(\Mux32~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~11 .lut_mask = 16'hBCB0;
defparam \Mux32~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y25_N19
dffeas \reg_file[2][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][31] .is_wysiwyg = "true";
defparam \reg_file[2][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N31
dffeas \reg_file[1][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][31] .is_wysiwyg = "true";
defparam \reg_file[1][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N21
dffeas \reg_file[3][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][31] .is_wysiwyg = "true";
defparam \reg_file[3][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N30
cycloneive_lcell_comb \Mux32~14 (
// Equation(s):
// \Mux32~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][31]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][31]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][31]~q ),
	.datad(\reg_file[3][31]~q ),
	.cin(gnd),
	.combout(\Mux32~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~14 .lut_mask = 16'hC840;
defparam \Mux32~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N18
cycloneive_lcell_comb \Mux32~15 (
// Equation(s):
// \Mux32~15_combout  = (\Mux32~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][31]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[2][31]~q ),
	.datad(\Mux32~14_combout ),
	.cin(gnd),
	.combout(\Mux32~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~15 .lut_mask = 16'hFF40;
defparam \Mux32~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y25_N1
dffeas \reg_file[10][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][31] .is_wysiwyg = "true";
defparam \reg_file[10][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N11
dffeas \reg_file[8][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][31] .is_wysiwyg = "true";
defparam \reg_file[8][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N10
cycloneive_lcell_comb \Mux32~12 (
// Equation(s):
// \Mux32~12_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[10][31]~q )) # (!\prif.imemload_id [17] & ((\reg_file[8][31]~q )))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[10][31]~q ),
	.datac(\reg_file[8][31]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux32~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~12 .lut_mask = 16'hEE50;
defparam \Mux32~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y25_N31
dffeas \reg_file[11][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][31] .is_wysiwyg = "true";
defparam \reg_file[11][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y25_N13
dffeas \reg_file[9][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][31] .is_wysiwyg = "true";
defparam \reg_file[9][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N30
cycloneive_lcell_comb \Mux32~13 (
// Equation(s):
// \Mux32~13_combout  = (\prif.imemload_id [16] & ((\Mux32~12_combout  & (\reg_file[11][31]~q )) # (!\Mux32~12_combout  & ((\reg_file[9][31]~q ))))) # (!\prif.imemload_id [16] & (\Mux32~12_combout ))

	.dataa(prifimemload_id_16),
	.datab(\Mux32~12_combout ),
	.datac(\reg_file[11][31]~q ),
	.datad(\reg_file[9][31]~q ),
	.cin(gnd),
	.combout(\Mux32~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~13 .lut_mask = 16'hE6C4;
defparam \Mux32~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N28
cycloneive_lcell_comb \Mux32~16 (
// Equation(s):
// \Mux32~16_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\Mux32~13_combout ))) # (!\prif.imemload_id [19] & (\Mux32~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux32~15_combout ),
	.datac(prifimemload_id_19),
	.datad(\Mux32~13_combout ),
	.cin(gnd),
	.combout(\Mux32~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux32~16 .lut_mask = 16'hF4A4;
defparam \Mux32~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N14
cycloneive_lcell_comb \reg_file_nxt[31][30]~70 (
// Equation(s):
// \reg_file_nxt[31][30]~70_combout  = (\Mux134~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Equal8),
	.datac(prifregwrite_wb_0),
	.datad(Mux134),
	.cin(gnd),
	.combout(\reg_file_nxt[31][30]~70_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][30]~70 .lut_mask = 16'hFB00;
defparam \reg_file_nxt[31][30]~70 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y27_N11
dffeas \reg_file[31][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][30] .is_wysiwyg = "true";
defparam \reg_file[31][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N5
dffeas \reg_file[27][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][30] .is_wysiwyg = "true";
defparam \reg_file[27][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N5
dffeas \reg_file[23][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][30] .is_wysiwyg = "true";
defparam \reg_file[23][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N23
dffeas \reg_file[19][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][30] .is_wysiwyg = "true";
defparam \reg_file[19][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N4
cycloneive_lcell_comb \Mux33~7 (
// Equation(s):
// \Mux33~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][30]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][30]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][30]~q ),
	.datad(\reg_file[19][30]~q ),
	.cin(gnd),
	.combout(\Mux33~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~7 .lut_mask = 16'hB9A8;
defparam \Mux33~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N4
cycloneive_lcell_comb \Mux33~8 (
// Equation(s):
// \Mux33~8_combout  = (\prif.imemload_id [19] & ((\Mux33~7_combout  & (\reg_file[31][30]~q )) # (!\Mux33~7_combout  & ((\reg_file[27][30]~q ))))) # (!\prif.imemload_id [19] & (((\Mux33~7_combout ))))

	.dataa(\reg_file[31][30]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][30]~q ),
	.datad(\Mux33~7_combout ),
	.cin(gnd),
	.combout(\Mux33~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~8 .lut_mask = 16'hBBC0;
defparam \Mux33~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N9
dffeas \reg_file[25][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][30] .is_wysiwyg = "true";
defparam \reg_file[25][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y27_N19
dffeas \reg_file[29][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][30] .is_wysiwyg = "true";
defparam \reg_file[29][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N7
dffeas \reg_file[17][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][30] .is_wysiwyg = "true";
defparam \reg_file[17][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N24
cycloneive_lcell_comb \reg_file[21][30]~feeder (
// Equation(s):
// \reg_file[21][30]~feeder_combout  = \reg_file_nxt[31][30]~70_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][30]~70_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[21][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][30]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[21][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N25
dffeas \reg_file[21][30] (
	.clk(!CLK),
	.d(\reg_file[21][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][30] .is_wysiwyg = "true";
defparam \reg_file[21][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N6
cycloneive_lcell_comb \Mux33~0 (
// Equation(s):
// \Mux33~0_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[21][30]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & (\reg_file[17][30]~q )))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][30]~q ),
	.datad(\reg_file[21][30]~q ),
	.cin(gnd),
	.combout(\Mux33~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~0 .lut_mask = 16'hBA98;
defparam \Mux33~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N18
cycloneive_lcell_comb \Mux33~1 (
// Equation(s):
// \Mux33~1_combout  = (\prif.imemload_id [19] & ((\Mux33~0_combout  & ((\reg_file[29][30]~q ))) # (!\Mux33~0_combout  & (\reg_file[25][30]~q )))) # (!\prif.imemload_id [19] & (((\Mux33~0_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[25][30]~q ),
	.datac(\reg_file[29][30]~q ),
	.datad(\Mux33~0_combout ),
	.cin(gnd),
	.combout(\Mux33~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~1 .lut_mask = 16'hF588;
defparam \Mux33~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y30_N13
dffeas \reg_file[18][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][30] .is_wysiwyg = "true";
defparam \reg_file[18][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N7
dffeas \reg_file[26][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][30] .is_wysiwyg = "true";
defparam \reg_file[26][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N12
cycloneive_lcell_comb \Mux33~2 (
// Equation(s):
// \Mux33~2_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[26][30]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & (\reg_file[18][30]~q )))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][30]~q ),
	.datad(\reg_file[26][30]~q ),
	.cin(gnd),
	.combout(\Mux33~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~2 .lut_mask = 16'hBA98;
defparam \Mux33~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N31
dffeas \reg_file[30][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][30] .is_wysiwyg = "true";
defparam \reg_file[30][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N25
dffeas \reg_file[22][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][30] .is_wysiwyg = "true";
defparam \reg_file[22][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N30
cycloneive_lcell_comb \Mux33~3 (
// Equation(s):
// \Mux33~3_combout  = (\prif.imemload_id [18] & ((\Mux33~2_combout  & (\reg_file[30][30]~q )) # (!\Mux33~2_combout  & ((\reg_file[22][30]~q ))))) # (!\prif.imemload_id [18] & (\Mux33~2_combout ))

	.dataa(prifimemload_id_18),
	.datab(\Mux33~2_combout ),
	.datac(\reg_file[30][30]~q ),
	.datad(\reg_file[22][30]~q ),
	.cin(gnd),
	.combout(\Mux33~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~3 .lut_mask = 16'hE6C4;
defparam \Mux33~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N20
cycloneive_lcell_comb \reg_file[28][30]~feeder (
// Equation(s):
// \reg_file[28][30]~feeder_combout  = \reg_file_nxt[31][30]~70_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][30]~70_combout ),
	.cin(gnd),
	.combout(\reg_file[28][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[28][30]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[28][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N21
dffeas \reg_file[28][30] (
	.clk(!CLK),
	.d(\reg_file[28][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][30] .is_wysiwyg = "true";
defparam \reg_file[28][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N17
dffeas \reg_file[20][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][30] .is_wysiwyg = "true";
defparam \reg_file[20][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N16
cycloneive_lcell_comb \Mux33~5 (
// Equation(s):
// \Mux33~5_combout  = (\Mux33~4_combout  & ((\reg_file[28][30]~q ) # ((!\prif.imemload_id [18])))) # (!\Mux33~4_combout  & (((\reg_file[20][30]~q  & \prif.imemload_id [18]))))

	.dataa(\Mux33~4_combout ),
	.datab(\reg_file[28][30]~q ),
	.datac(\reg_file[20][30]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux33~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~5 .lut_mask = 16'hD8AA;
defparam \Mux33~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N12
cycloneive_lcell_comb \Mux33~6 (
// Equation(s):
// \Mux33~6_combout  = (\prif.imemload_id [17] & ((\Mux33~3_combout ) # ((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (((!\prif.imemload_id [16] & \Mux33~5_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\Mux33~3_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux33~5_combout ),
	.cin(gnd),
	.combout(\Mux33~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~6 .lut_mask = 16'hADA8;
defparam \Mux33~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N17
dffeas \reg_file[6][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][30] .is_wysiwyg = "true";
defparam \reg_file[6][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N9
dffeas \reg_file[5][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][30] .is_wysiwyg = "true";
defparam \reg_file[5][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N3
dffeas \reg_file[4][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][30] .is_wysiwyg = "true";
defparam \reg_file[4][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N2
cycloneive_lcell_comb \Mux33~12 (
// Equation(s):
// \Mux33~12_combout  = (\prif.imemload_id [16] & ((\reg_file[5][30]~q ) # ((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & (((\reg_file[4][30]~q  & !\prif.imemload_id [17]))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[5][30]~q ),
	.datac(\reg_file[4][30]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux33~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~12 .lut_mask = 16'hAAD8;
defparam \Mux33~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N18
cycloneive_lcell_comb \Mux33~13 (
// Equation(s):
// \Mux33~13_combout  = (\Mux33~12_combout  & ((\reg_file[7][30]~q ) # ((!\prif.imemload_id [17])))) # (!\Mux33~12_combout  & (((\reg_file[6][30]~q  & \prif.imemload_id [17]))))

	.dataa(\reg_file[7][30]~q ),
	.datab(\reg_file[6][30]~q ),
	.datac(\Mux33~12_combout ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux33~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~13 .lut_mask = 16'hACF0;
defparam \Mux33~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N21
dffeas \reg_file[2][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][30] .is_wysiwyg = "true";
defparam \reg_file[2][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N20
cycloneive_lcell_comb \Mux33~15 (
// Equation(s):
// \Mux33~15_combout  = (\Mux33~14_combout ) # ((!\prif.imemload_id [16] & (\reg_file[2][30]~q  & \prif.imemload_id [17])))

	.dataa(\Mux33~14_combout ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[2][30]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux33~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~15 .lut_mask = 16'hBAAA;
defparam \Mux33~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N30
cycloneive_lcell_comb \Mux33~16 (
// Equation(s):
// \Mux33~16_combout  = (\prif.imemload_id [18] & ((\Mux33~13_combout ) # ((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (((!\prif.imemload_id [19] & \Mux33~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux33~13_combout ),
	.datac(prifimemload_id_19),
	.datad(\Mux33~15_combout ),
	.cin(gnd),
	.combout(\Mux33~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~16 .lut_mask = 16'hADA8;
defparam \Mux33~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N15
dffeas \reg_file[14][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][30] .is_wysiwyg = "true";
defparam \reg_file[14][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N11
dffeas \reg_file[12][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][30] .is_wysiwyg = "true";
defparam \reg_file[12][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N13
dffeas \reg_file[13][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][30] .is_wysiwyg = "true";
defparam \reg_file[13][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N10
cycloneive_lcell_comb \Mux33~17 (
// Equation(s):
// \Mux33~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][30]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][30]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][30]~q ),
	.datad(\reg_file[13][30]~q ),
	.cin(gnd),
	.combout(\Mux33~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~17 .lut_mask = 16'hDC98;
defparam \Mux33~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N15
dffeas \reg_file[15][30] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][30]~70_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][30] .is_wysiwyg = "true";
defparam \reg_file[15][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N8
cycloneive_lcell_comb \Mux33~18 (
// Equation(s):
// \Mux33~18_combout  = (\prif.imemload_id [17] & ((\Mux33~17_combout  & ((\reg_file[15][30]~q ))) # (!\Mux33~17_combout  & (\reg_file[14][30]~q )))) # (!\prif.imemload_id [17] & (((\Mux33~17_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[14][30]~q ),
	.datac(\Mux33~17_combout ),
	.datad(\reg_file[15][30]~q ),
	.cin(gnd),
	.combout(\Mux33~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~18 .lut_mask = 16'hF858;
defparam \Mux33~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y25_N19
dffeas \reg_file[11][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][30] .is_wysiwyg = "true";
defparam \reg_file[11][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y25_N21
dffeas \reg_file[9][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][30] .is_wysiwyg = "true";
defparam \reg_file[9][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N15
dffeas \reg_file[8][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][30] .is_wysiwyg = "true";
defparam \reg_file[8][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N25
dffeas \reg_file[10][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][30] .is_wysiwyg = "true";
defparam \reg_file[10][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N24
cycloneive_lcell_comb \Mux33~10 (
// Equation(s):
// \Mux33~10_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][30]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][30]~q ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[8][30]~q ),
	.datac(\reg_file[10][30]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux33~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~10 .lut_mask = 16'hFA44;
defparam \Mux33~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N20
cycloneive_lcell_comb \Mux33~11 (
// Equation(s):
// \Mux33~11_combout  = (\prif.imemload_id [16] & ((\Mux33~10_combout  & (\reg_file[11][30]~q )) # (!\Mux33~10_combout  & ((\reg_file[9][30]~q ))))) # (!\prif.imemload_id [16] & (((\Mux33~10_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[11][30]~q ),
	.datac(\reg_file[9][30]~q ),
	.datad(\Mux33~10_combout ),
	.cin(gnd),
	.combout(\Mux33~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux33~11 .lut_mask = 16'hDDA0;
defparam \Mux33~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N6
cycloneive_lcell_comb \reg_file_nxt[31][29]~71 (
// Equation(s):
// \reg_file_nxt[31][29]~71_combout  = (\Mux135~1_combout  & (((\prif.regwrite_wb [2]) # (\prif.regwrite_wb [0])) # (!Equal8)))

	.dataa(Equal8),
	.datab(prifregwrite_wb_2),
	.datac(Mux135),
	.datad(prifregwrite_wb_0),
	.cin(gnd),
	.combout(\reg_file_nxt[31][29]~71_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][29]~71 .lut_mask = 16'hF0D0;
defparam \reg_file_nxt[31][29]~71 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y26_N9
dffeas \reg_file[27][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][29] .is_wysiwyg = "true";
defparam \reg_file[27][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N25
dffeas \reg_file[19][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][29] .is_wysiwyg = "true";
defparam \reg_file[19][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N8
cycloneive_lcell_comb \Mux34~7 (
// Equation(s):
// \Mux34~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][29]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][29]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][29]~q ),
	.datad(\reg_file[19][29]~q ),
	.cin(gnd),
	.combout(\Mux34~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~7 .lut_mask = 16'hD9C8;
defparam \Mux34~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N11
dffeas \reg_file[23][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][29] .is_wysiwyg = "true";
defparam \reg_file[23][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y26_N19
dffeas \reg_file[31][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][29] .is_wysiwyg = "true";
defparam \reg_file[31][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N10
cycloneive_lcell_comb \Mux34~8 (
// Equation(s):
// \Mux34~8_combout  = (\prif.imemload_id [18] & ((\Mux34~7_combout  & ((\reg_file[31][29]~q ))) # (!\Mux34~7_combout  & (\reg_file[23][29]~q )))) # (!\prif.imemload_id [18] & (\Mux34~7_combout ))

	.dataa(prifimemload_id_18),
	.datab(\Mux34~7_combout ),
	.datac(\reg_file[23][29]~q ),
	.datad(\reg_file[31][29]~q ),
	.cin(gnd),
	.combout(\Mux34~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~8 .lut_mask = 16'hEC64;
defparam \Mux34~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N2
cycloneive_lcell_comb \reg_file[29][29]~feeder (
// Equation(s):
// \reg_file[29][29]~feeder_combout  = \reg_file_nxt[31][29]~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][29]~71_combout ),
	.cin(gnd),
	.combout(\reg_file[29][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][29]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N3
dffeas \reg_file[29][29] (
	.clk(!CLK),
	.d(\reg_file[29][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][29] .is_wysiwyg = "true";
defparam \reg_file[29][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N1
dffeas \reg_file[17][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][29] .is_wysiwyg = "true";
defparam \reg_file[17][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N16
cycloneive_lcell_comb \reg_file[25][29]~feeder (
// Equation(s):
// \reg_file[25][29]~feeder_combout  = \reg_file_nxt[31][29]~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][29]~71_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[25][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][29]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[25][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N17
dffeas \reg_file[25][29] (
	.clk(!CLK),
	.d(\reg_file[25][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][29] .is_wysiwyg = "true";
defparam \reg_file[25][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N0
cycloneive_lcell_comb \Mux34~0 (
// Equation(s):
// \Mux34~0_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[25][29]~q ))) # (!\prif.imemload_id [19] & (\reg_file[17][29]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][29]~q ),
	.datad(\reg_file[25][29]~q ),
	.cin(gnd),
	.combout(\Mux34~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~0 .lut_mask = 16'hDC98;
defparam \Mux34~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N31
dffeas \reg_file[21][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][29] .is_wysiwyg = "true";
defparam \reg_file[21][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N4
cycloneive_lcell_comb \Mux34~1 (
// Equation(s):
// \Mux34~1_combout  = (\prif.imemload_id [18] & ((\Mux34~0_combout  & (\reg_file[29][29]~q )) # (!\Mux34~0_combout  & ((\reg_file[21][29]~q ))))) # (!\prif.imemload_id [18] & (((\Mux34~0_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[29][29]~q ),
	.datac(\Mux34~0_combout ),
	.datad(\reg_file[21][29]~q ),
	.cin(gnd),
	.combout(\Mux34~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~1 .lut_mask = 16'hDAD0;
defparam \Mux34~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N21
dffeas \reg_file[26][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][29] .is_wysiwyg = "true";
defparam \reg_file[26][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N7
dffeas \reg_file[30][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][29] .is_wysiwyg = "true";
defparam \reg_file[30][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N19
dffeas \reg_file[18][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][29] .is_wysiwyg = "true";
defparam \reg_file[18][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N17
dffeas \reg_file[22][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][29] .is_wysiwyg = "true";
defparam \reg_file[22][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N18
cycloneive_lcell_comb \Mux34~2 (
// Equation(s):
// \Mux34~2_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[22][29]~q ))) # (!\prif.imemload_id [18] & (\reg_file[18][29]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][29]~q ),
	.datad(\reg_file[22][29]~q ),
	.cin(gnd),
	.combout(\Mux34~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~2 .lut_mask = 16'hDC98;
defparam \Mux34~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N6
cycloneive_lcell_comb \Mux34~3 (
// Equation(s):
// \Mux34~3_combout  = (\prif.imemload_id [19] & ((\Mux34~2_combout  & ((\reg_file[30][29]~q ))) # (!\Mux34~2_combout  & (\reg_file[26][29]~q )))) # (!\prif.imemload_id [19] & (((\Mux34~2_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[26][29]~q ),
	.datac(\reg_file[30][29]~q ),
	.datad(\Mux34~2_combout ),
	.cin(gnd),
	.combout(\Mux34~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~3 .lut_mask = 16'hF588;
defparam \Mux34~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N15
dffeas \reg_file[28][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][29] .is_wysiwyg = "true";
defparam \reg_file[28][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N21
dffeas \reg_file[24][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][29] .is_wysiwyg = "true";
defparam \reg_file[24][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N20
cycloneive_lcell_comb \Mux34~5 (
// Equation(s):
// \Mux34~5_combout  = (\Mux34~4_combout  & ((\reg_file[28][29]~q ) # ((!\prif.imemload_id [19])))) # (!\Mux34~4_combout  & (((\reg_file[24][29]~q  & \prif.imemload_id [19]))))

	.dataa(\Mux34~4_combout ),
	.datab(\reg_file[28][29]~q ),
	.datac(\reg_file[24][29]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux34~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~5 .lut_mask = 16'hD8AA;
defparam \Mux34~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N12
cycloneive_lcell_comb \Mux34~6 (
// Equation(s):
// \Mux34~6_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\Mux34~3_combout )) # (!\prif.imemload_id [17] & ((\Mux34~5_combout )))))

	.dataa(prifimemload_id_16),
	.datab(\Mux34~3_combout ),
	.datac(prifimemload_id_17),
	.datad(\Mux34~5_combout ),
	.cin(gnd),
	.combout(\Mux34~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~6 .lut_mask = 16'hE5E0;
defparam \Mux34~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N24
cycloneive_lcell_comb \reg_file[14][29]~feeder (
// Equation(s):
// \reg_file[14][29]~feeder_combout  = \reg_file_nxt[31][29]~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][29]~71_combout ),
	.cin(gnd),
	.combout(\reg_file[14][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][29]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[14][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N25
dffeas \reg_file[14][29] (
	.clk(!CLK),
	.d(\reg_file[14][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][29] .is_wysiwyg = "true";
defparam \reg_file[14][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N3
dffeas \reg_file[12][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][29] .is_wysiwyg = "true";
defparam \reg_file[12][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N21
dffeas \reg_file[13][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][29] .is_wysiwyg = "true";
defparam \reg_file[13][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N2
cycloneive_lcell_comb \Mux34~17 (
// Equation(s):
// \Mux34~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][29]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][29]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][29]~q ),
	.datad(\reg_file[13][29]~q ),
	.cin(gnd),
	.combout(\Mux34~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~17 .lut_mask = 16'hDC98;
defparam \Mux34~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N28
cycloneive_lcell_comb \reg_file[15][29]~feeder (
// Equation(s):
// \reg_file[15][29]~feeder_combout  = \reg_file_nxt[31][29]~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][29]~71_combout ),
	.cin(gnd),
	.combout(\reg_file[15][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[15][29]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[15][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N29
dffeas \reg_file[15][29] (
	.clk(!CLK),
	.d(\reg_file[15][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][29] .is_wysiwyg = "true";
defparam \reg_file[15][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N0
cycloneive_lcell_comb \Mux34~18 (
// Equation(s):
// \Mux34~18_combout  = (\Mux34~17_combout  & (((\reg_file[15][29]~q ) # (!\prif.imemload_id [17])))) # (!\Mux34~17_combout  & (\reg_file[14][29]~q  & ((\prif.imemload_id [17]))))

	.dataa(\reg_file[14][29]~q ),
	.datab(\Mux34~17_combout ),
	.datac(\reg_file[15][29]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux34~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~18 .lut_mask = 16'hE2CC;
defparam \Mux34~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N5
dffeas \reg_file[2][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][29] .is_wysiwyg = "true";
defparam \reg_file[2][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N25
dffeas \reg_file[1][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][29] .is_wysiwyg = "true";
defparam \reg_file[1][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N15
dffeas \reg_file[3][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][29] .is_wysiwyg = "true";
defparam \reg_file[3][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N24
cycloneive_lcell_comb \Mux34~14 (
// Equation(s):
// \Mux34~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][29]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][29]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][29]~q ),
	.datad(\reg_file[3][29]~q ),
	.cin(gnd),
	.combout(\Mux34~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~14 .lut_mask = 16'hC840;
defparam \Mux34~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N4
cycloneive_lcell_comb \Mux34~15 (
// Equation(s):
// \Mux34~15_combout  = (\Mux34~14_combout ) # ((\prif.imemload_id [17] & (!\prif.imemload_id [16] & \reg_file[2][29]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[2][29]~q ),
	.datad(\Mux34~14_combout ),
	.cin(gnd),
	.combout(\Mux34~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~15 .lut_mask = 16'hFF20;
defparam \Mux34~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N7
dffeas \reg_file[11][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][29] .is_wysiwyg = "true";
defparam \reg_file[11][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N1
dffeas \reg_file[10][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][29] .is_wysiwyg = "true";
defparam \reg_file[10][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N19
dffeas \reg_file[8][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][29] .is_wysiwyg = "true";
defparam \reg_file[8][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N0
cycloneive_lcell_comb \Mux34~12 (
// Equation(s):
// \Mux34~12_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[10][29]~q )) # (!\prif.imemload_id [17] & ((\reg_file[8][29]~q )))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[10][29]~q ),
	.datad(\reg_file[8][29]~q ),
	.cin(gnd),
	.combout(\Mux34~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~12 .lut_mask = 16'hD9C8;
defparam \Mux34~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N6
cycloneive_lcell_comb \Mux34~13 (
// Equation(s):
// \Mux34~13_combout  = (\prif.imemload_id [16] & ((\Mux34~12_combout  & ((\reg_file[11][29]~q ))) # (!\Mux34~12_combout  & (\reg_file[9][29]~q )))) # (!\prif.imemload_id [16] & (((\Mux34~12_combout ))))

	.dataa(\reg_file[9][29]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[11][29]~q ),
	.datad(\Mux34~12_combout ),
	.cin(gnd),
	.combout(\Mux34~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~13 .lut_mask = 16'hF388;
defparam \Mux34~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N22
cycloneive_lcell_comb \Mux34~16 (
// Equation(s):
// \Mux34~16_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\Mux34~13_combout ))) # (!\prif.imemload_id [19] & (\Mux34~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\Mux34~15_combout ),
	.datac(prifimemload_id_19),
	.datad(\Mux34~13_combout ),
	.cin(gnd),
	.combout(\Mux34~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~16 .lut_mask = 16'hF4A4;
defparam \Mux34~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N17
dffeas \reg_file[4][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][29] .is_wysiwyg = "true";
defparam \reg_file[4][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N27
dffeas \reg_file[5][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][29] .is_wysiwyg = "true";
defparam \reg_file[5][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N26
cycloneive_lcell_comb \Mux34~10 (
// Equation(s):
// \Mux34~10_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[5][29]~q ))) # (!\prif.imemload_id [16] & (\reg_file[4][29]~q ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[4][29]~q ),
	.datac(\reg_file[5][29]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux34~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~10 .lut_mask = 16'hFA44;
defparam \Mux34~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N25
dffeas \reg_file[6][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][29] .is_wysiwyg = "true";
defparam \reg_file[6][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N11
dffeas \reg_file[7][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][29] .is_wysiwyg = "true";
defparam \reg_file[7][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N24
cycloneive_lcell_comb \Mux34~11 (
// Equation(s):
// \Mux34~11_combout  = (\prif.imemload_id [17] & ((\Mux34~10_combout  & ((\reg_file[7][29]~q ))) # (!\Mux34~10_combout  & (\reg_file[6][29]~q )))) # (!\prif.imemload_id [17] & (\Mux34~10_combout ))

	.dataa(prifimemload_id_17),
	.datab(\Mux34~10_combout ),
	.datac(\reg_file[6][29]~q ),
	.datad(\reg_file[7][29]~q ),
	.cin(gnd),
	.combout(\Mux34~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux34~11 .lut_mask = 16'hEC64;
defparam \Mux34~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N28
cycloneive_lcell_comb \reg_file_nxt[31][5]~72 (
// Equation(s):
// \reg_file_nxt[31][5]~72_combout  = (\Mux159~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Mux159),
	.datac(prifregwrite_wb_0),
	.datad(Equal8),
	.cin(gnd),
	.combout(\reg_file_nxt[31][5]~72_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][5]~72 .lut_mask = 16'hC8CC;
defparam \reg_file_nxt[31][5]~72 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N27
dffeas \reg_file[30][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][5] .is_wysiwyg = "true";
defparam \reg_file[30][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N15
dffeas \reg_file[26][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][5] .is_wysiwyg = "true";
defparam \reg_file[26][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N8
cycloneive_lcell_comb \Mux58~3 (
// Equation(s):
// \Mux58~3_combout  = (\Mux58~2_combout  & ((\reg_file[30][5]~q ) # ((!\prif.imemload_id [19])))) # (!\Mux58~2_combout  & (((\reg_file[26][5]~q  & \prif.imemload_id [19]))))

	.dataa(\Mux58~2_combout ),
	.datab(\reg_file[30][5]~q ),
	.datac(\reg_file[26][5]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux58~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~3 .lut_mask = 16'hD8AA;
defparam \Mux58~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N17
dffeas \reg_file[24][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][5] .is_wysiwyg = "true";
defparam \reg_file[24][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N9
dffeas \reg_file[20][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][5] .is_wysiwyg = "true";
defparam \reg_file[20][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N19
dffeas \reg_file[16][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][5] .is_wysiwyg = "true";
defparam \reg_file[16][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N8
cycloneive_lcell_comb \Mux58~4 (
// Equation(s):
// \Mux58~4_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[20][5]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[16][5]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[20][5]~q ),
	.datad(\reg_file[16][5]~q ),
	.cin(gnd),
	.combout(\Mux58~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~4 .lut_mask = 16'hB9A8;
defparam \Mux58~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N16
cycloneive_lcell_comb \Mux58~5 (
// Equation(s):
// \Mux58~5_combout  = (\prif.imemload_id [19] & ((\Mux58~4_combout  & (\reg_file[28][5]~q )) # (!\Mux58~4_combout  & ((\reg_file[24][5]~q ))))) # (!\prif.imemload_id [19] & (((\Mux58~4_combout ))))

	.dataa(\reg_file[28][5]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[24][5]~q ),
	.datad(\Mux58~4_combout ),
	.cin(gnd),
	.combout(\Mux58~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~5 .lut_mask = 16'hBBC0;
defparam \Mux58~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N18
cycloneive_lcell_comb \Mux58~6 (
// Equation(s):
// \Mux58~6_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\Mux58~3_combout )) # (!\prif.imemload_id [17] & ((\Mux58~5_combout )))))

	.dataa(prifimemload_id_16),
	.datab(\Mux58~3_combout ),
	.datac(prifimemload_id_17),
	.datad(\Mux58~5_combout ),
	.cin(gnd),
	.combout(\Mux58~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~6 .lut_mask = 16'hE5E0;
defparam \Mux58~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N13
dffeas \reg_file[25][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][5] .is_wysiwyg = "true";
defparam \reg_file[25][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y26_N5
dffeas \reg_file[17][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][5] .is_wysiwyg = "true";
defparam \reg_file[17][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N12
cycloneive_lcell_comb \Mux58~0 (
// Equation(s):
// \Mux58~0_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[25][5]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & ((\reg_file[17][5]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[25][5]~q ),
	.datad(\reg_file[17][5]~q ),
	.cin(gnd),
	.combout(\Mux58~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~0 .lut_mask = 16'hB9A8;
defparam \Mux58~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N12
cycloneive_lcell_comb \reg_file[21][5]~feeder (
// Equation(s):
// \reg_file[21][5]~feeder_combout  = \reg_file_nxt[31][5]~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][5]~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[21][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][5]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[21][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N13
dffeas \reg_file[21][5] (
	.clk(!CLK),
	.d(\reg_file[21][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][5] .is_wysiwyg = "true";
defparam \reg_file[21][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N14
cycloneive_lcell_comb \reg_file[29][5]~feeder (
// Equation(s):
// \reg_file[29][5]~feeder_combout  = \reg_file_nxt[31][5]~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][5]~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][5]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N15
dffeas \reg_file[29][5] (
	.clk(!CLK),
	.d(\reg_file[29][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][5] .is_wysiwyg = "true";
defparam \reg_file[29][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N10
cycloneive_lcell_comb \Mux58~1 (
// Equation(s):
// \Mux58~1_combout  = (\prif.imemload_id [18] & ((\Mux58~0_combout  & ((\reg_file[29][5]~q ))) # (!\Mux58~0_combout  & (\reg_file[21][5]~q )))) # (!\prif.imemload_id [18] & (\Mux58~0_combout ))

	.dataa(prifimemload_id_18),
	.datab(\Mux58~0_combout ),
	.datac(\reg_file[21][5]~q ),
	.datad(\reg_file[29][5]~q ),
	.cin(gnd),
	.combout(\Mux58~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~1 .lut_mask = 16'hEC64;
defparam \Mux58~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N10
cycloneive_lcell_comb \reg_file[23][5]~feeder (
// Equation(s):
// \reg_file[23][5]~feeder_combout  = \reg_file_nxt[31][5]~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][5]~72_combout ),
	.cin(gnd),
	.combout(\reg_file[23][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][5]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[23][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N11
dffeas \reg_file[23][5] (
	.clk(!CLK),
	.d(\reg_file[23][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][5] .is_wysiwyg = "true";
defparam \reg_file[23][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N24
cycloneive_lcell_comb \reg_file[31][5]~feeder (
// Equation(s):
// \reg_file[31][5]~feeder_combout  = \reg_file_nxt[31][5]~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][5]~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[31][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][5]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[31][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y26_N25
dffeas \reg_file[31][5] (
	.clk(!CLK),
	.d(\reg_file[31][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][5] .is_wysiwyg = "true";
defparam \reg_file[31][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y26_N29
dffeas \reg_file[27][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][5] .is_wysiwyg = "true";
defparam \reg_file[27][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N3
dffeas \reg_file[19][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][5] .is_wysiwyg = "true";
defparam \reg_file[19][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N28
cycloneive_lcell_comb \Mux58~7 (
// Equation(s):
// \Mux58~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][5]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][5]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][5]~q ),
	.datad(\reg_file[19][5]~q ),
	.cin(gnd),
	.combout(\Mux58~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~7 .lut_mask = 16'hD9C8;
defparam \Mux58~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N18
cycloneive_lcell_comb \Mux58~8 (
// Equation(s):
// \Mux58~8_combout  = (\prif.imemload_id [18] & ((\Mux58~7_combout  & ((\reg_file[31][5]~q ))) # (!\Mux58~7_combout  & (\reg_file[23][5]~q )))) # (!\prif.imemload_id [18] & (((\Mux58~7_combout ))))

	.dataa(\reg_file[23][5]~q ),
	.datab(\reg_file[31][5]~q ),
	.datac(prifimemload_id_18),
	.datad(\Mux58~7_combout ),
	.cin(gnd),
	.combout(\Mux58~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~8 .lut_mask = 16'hCFA0;
defparam \Mux58~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N24
cycloneive_lcell_comb \reg_file[6][5]~feeder (
// Equation(s):
// \reg_file[6][5]~feeder_combout  = \reg_file_nxt[31][5]~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][5]~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][5]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N25
dffeas \reg_file[6][5] (
	.clk(!CLK),
	.d(\reg_file[6][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][5] .is_wysiwyg = "true";
defparam \reg_file[6][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N31
dffeas \reg_file[7][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][5] .is_wysiwyg = "true";
defparam \reg_file[7][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N5
dffeas \reg_file[4][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][5] .is_wysiwyg = "true";
defparam \reg_file[4][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N21
dffeas \reg_file[5][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][5] .is_wysiwyg = "true";
defparam \reg_file[5][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N20
cycloneive_lcell_comb \Mux58~10 (
// Equation(s):
// \Mux58~10_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[5][5]~q ))) # (!\prif.imemload_id [16] & (\reg_file[4][5]~q ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[4][5]~q ),
	.datac(\reg_file[5][5]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux58~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~10 .lut_mask = 16'hFA44;
defparam \Mux58~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N26
cycloneive_lcell_comb \Mux58~11 (
// Equation(s):
// \Mux58~11_combout  = (\prif.imemload_id [17] & ((\Mux58~10_combout  & ((\reg_file[7][5]~q ))) # (!\Mux58~10_combout  & (\reg_file[6][5]~q )))) # (!\prif.imemload_id [17] & (((\Mux58~10_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][5]~q ),
	.datac(\reg_file[7][5]~q ),
	.datad(\Mux58~10_combout ),
	.cin(gnd),
	.combout(\Mux58~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~11 .lut_mask = 16'hF588;
defparam \Mux58~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y27_N1
dffeas \reg_file[1][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][5] .is_wysiwyg = "true";
defparam \reg_file[1][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N3
dffeas \reg_file[3][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][5] .is_wysiwyg = "true";
defparam \reg_file[3][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N0
cycloneive_lcell_comb \Mux58~14 (
// Equation(s):
// \Mux58~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][5]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][5]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][5]~q ),
	.datad(\reg_file[3][5]~q ),
	.cin(gnd),
	.combout(\Mux58~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~14 .lut_mask = 16'hC840;
defparam \Mux58~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N12
cycloneive_lcell_comb \Mux58~15 (
// Equation(s):
// \Mux58~15_combout  = (\Mux58~14_combout ) # ((\reg_file[2][5]~q  & (\prif.imemload_id [17] & !\prif.imemload_id [16])))

	.dataa(\reg_file[2][5]~q ),
	.datab(\Mux58~14_combout ),
	.datac(prifimemload_id_17),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux58~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~15 .lut_mask = 16'hCCEC;
defparam \Mux58~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N22
cycloneive_lcell_comb \reg_file[9][5]~feeder (
// Equation(s):
// \reg_file[9][5]~feeder_combout  = \reg_file_nxt[31][5]~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][5]~72_combout ),
	.cin(gnd),
	.combout(\reg_file[9][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[9][5]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[9][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N23
dffeas \reg_file[9][5] (
	.clk(!CLK),
	.d(\reg_file[9][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][5] .is_wysiwyg = "true";
defparam \reg_file[9][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N21
dffeas \reg_file[11][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][5] .is_wysiwyg = "true";
defparam \reg_file[11][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N5
dffeas \reg_file[10][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][5] .is_wysiwyg = "true";
defparam \reg_file[10][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N3
dffeas \reg_file[8][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][5] .is_wysiwyg = "true";
defparam \reg_file[8][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N2
cycloneive_lcell_comb \Mux58~12 (
// Equation(s):
// \Mux58~12_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[10][5]~q )) # (!\prif.imemload_id [17] & ((\reg_file[8][5]~q )))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[10][5]~q ),
	.datac(\reg_file[8][5]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux58~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~12 .lut_mask = 16'hEE50;
defparam \Mux58~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N20
cycloneive_lcell_comb \Mux58~13 (
// Equation(s):
// \Mux58~13_combout  = (\prif.imemload_id [16] & ((\Mux58~12_combout  & ((\reg_file[11][5]~q ))) # (!\Mux58~12_combout  & (\reg_file[9][5]~q )))) # (!\prif.imemload_id [16] & (((\Mux58~12_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[9][5]~q ),
	.datac(\reg_file[11][5]~q ),
	.datad(\Mux58~12_combout ),
	.cin(gnd),
	.combout(\Mux58~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~13 .lut_mask = 16'hF588;
defparam \Mux58~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N22
cycloneive_lcell_comb \Mux58~16 (
// Equation(s):
// \Mux58~16_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\Mux58~13_combout ))) # (!\prif.imemload_id [19] & (\Mux58~15_combout ))))

	.dataa(\Mux58~15_combout ),
	.datab(\Mux58~13_combout ),
	.datac(prifimemload_id_18),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux58~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~16 .lut_mask = 16'hFC0A;
defparam \Mux58~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y26_N9
dffeas \reg_file[13][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][5] .is_wysiwyg = "true";
defparam \reg_file[13][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N23
dffeas \reg_file[12][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][5] .is_wysiwyg = "true";
defparam \reg_file[12][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N22
cycloneive_lcell_comb \Mux58~17 (
// Equation(s):
// \Mux58~17_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & (\reg_file[13][5]~q )) # (!\prif.imemload_id [16] & ((\reg_file[12][5]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[13][5]~q ),
	.datac(\reg_file[12][5]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux58~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~17 .lut_mask = 16'hEE50;
defparam \Mux58~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N4
cycloneive_lcell_comb \reg_file[14][5]~feeder (
// Equation(s):
// \reg_file[14][5]~feeder_combout  = \reg_file_nxt[31][5]~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][5]~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[14][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][5]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[14][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y28_N5
dffeas \reg_file[14][5] (
	.clk(!CLK),
	.d(\reg_file[14][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][5] .is_wysiwyg = "true";
defparam \reg_file[14][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N29
dffeas \reg_file[15][5] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][5]~72_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][5] .is_wysiwyg = "true";
defparam \reg_file[15][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N2
cycloneive_lcell_comb \Mux58~18 (
// Equation(s):
// \Mux58~18_combout  = (\Mux58~17_combout  & (((\reg_file[15][5]~q ) # (!\prif.imemload_id [17])))) # (!\Mux58~17_combout  & (\reg_file[14][5]~q  & ((\prif.imemload_id [17]))))

	.dataa(\Mux58~17_combout ),
	.datab(\reg_file[14][5]~q ),
	.datac(\reg_file[15][5]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux58~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux58~18 .lut_mask = 16'hE4AA;
defparam \Mux58~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N26
cycloneive_lcell_comb \reg_file_nxt[31][15]~73 (
// Equation(s):
// \reg_file_nxt[31][15]~73_combout  = (\Mux149~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Equal8),
	.datac(prifregwrite_wb_0),
	.datad(Mux149),
	.cin(gnd),
	.combout(\reg_file_nxt[31][15]~73_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][15]~73 .lut_mask = 16'hFB00;
defparam \reg_file_nxt[31][15]~73 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N8
cycloneive_lcell_comb \reg_file[29][15]~feeder (
// Equation(s):
// \reg_file[29][15]~feeder_combout  = \reg_file_nxt[31][15]~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][15]~73_combout ),
	.cin(gnd),
	.combout(\reg_file[29][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][15]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N9
dffeas \reg_file[29][15] (
	.clk(!CLK),
	.d(\reg_file[29][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][15] .is_wysiwyg = "true";
defparam \reg_file[29][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y26_N5
dffeas \reg_file[21][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][15] .is_wysiwyg = "true";
defparam \reg_file[21][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y26_N19
dffeas \reg_file[17][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][15] .is_wysiwyg = "true";
defparam \reg_file[17][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y26_N7
dffeas \reg_file[25][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][15] .is_wysiwyg = "true";
defparam \reg_file[25][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N6
cycloneive_lcell_comb \Mux48~0 (
// Equation(s):
// \Mux48~0_combout  = (\prif.imemload_id [19] & (((\reg_file[25][15]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[17][15]~q  & ((!\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[17][15]~q ),
	.datac(\reg_file[25][15]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux48~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~0 .lut_mask = 16'hAAE4;
defparam \Mux48~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N4
cycloneive_lcell_comb \Mux48~1 (
// Equation(s):
// \Mux48~1_combout  = (\prif.imemload_id [18] & ((\Mux48~0_combout  & (\reg_file[29][15]~q )) # (!\Mux48~0_combout  & ((\reg_file[21][15]~q ))))) # (!\prif.imemload_id [18] & (((\Mux48~0_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[29][15]~q ),
	.datac(\reg_file[21][15]~q ),
	.datad(\Mux48~0_combout ),
	.cin(gnd),
	.combout(\Mux48~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~1 .lut_mask = 16'hDDA0;
defparam \Mux48~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y26_N3
dffeas \reg_file[27][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][15] .is_wysiwyg = "true";
defparam \reg_file[27][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N13
dffeas \reg_file[19][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][15] .is_wysiwyg = "true";
defparam \reg_file[19][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N2
cycloneive_lcell_comb \Mux48~7 (
// Equation(s):
// \Mux48~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][15]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][15]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][15]~q ),
	.datad(\reg_file[19][15]~q ),
	.cin(gnd),
	.combout(\Mux48~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~7 .lut_mask = 16'hD9C8;
defparam \Mux48~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y26_N13
dffeas \reg_file[31][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][15] .is_wysiwyg = "true";
defparam \reg_file[31][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N18
cycloneive_lcell_comb \reg_file[23][15]~feeder (
// Equation(s):
// \reg_file[23][15]~feeder_combout  = \reg_file_nxt[31][15]~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][15]~73_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[23][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][15]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[23][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y26_N19
dffeas \reg_file[23][15] (
	.clk(!CLK),
	.d(\reg_file[23][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][15] .is_wysiwyg = "true";
defparam \reg_file[23][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N12
cycloneive_lcell_comb \Mux48~8 (
// Equation(s):
// \Mux48~8_combout  = (\prif.imemload_id [18] & ((\Mux48~7_combout  & (\reg_file[31][15]~q )) # (!\Mux48~7_combout  & ((\reg_file[23][15]~q ))))) # (!\prif.imemload_id [18] & (\Mux48~7_combout ))

	.dataa(prifimemload_id_18),
	.datab(\Mux48~7_combout ),
	.datac(\reg_file[31][15]~q ),
	.datad(\reg_file[23][15]~q ),
	.cin(gnd),
	.combout(\Mux48~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~8 .lut_mask = 16'hE6C4;
defparam \Mux48~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N5
dffeas \reg_file[28][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][15] .is_wysiwyg = "true";
defparam \reg_file[28][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N15
dffeas \reg_file[24][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][15] .is_wysiwyg = "true";
defparam \reg_file[24][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N5
dffeas \reg_file[20][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][15] .is_wysiwyg = "true";
defparam \reg_file[20][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N11
dffeas \reg_file[16][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][15] .is_wysiwyg = "true";
defparam \reg_file[16][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N4
cycloneive_lcell_comb \Mux48~4 (
// Equation(s):
// \Mux48~4_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[20][15]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[16][15]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[20][15]~q ),
	.datad(\reg_file[16][15]~q ),
	.cin(gnd),
	.combout(\Mux48~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~4 .lut_mask = 16'hB9A8;
defparam \Mux48~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N14
cycloneive_lcell_comb \Mux48~5 (
// Equation(s):
// \Mux48~5_combout  = (\prif.imemload_id [19] & ((\Mux48~4_combout  & (\reg_file[28][15]~q )) # (!\Mux48~4_combout  & ((\reg_file[24][15]~q ))))) # (!\prif.imemload_id [19] & (((\Mux48~4_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[28][15]~q ),
	.datac(\reg_file[24][15]~q ),
	.datad(\Mux48~4_combout ),
	.cin(gnd),
	.combout(\Mux48~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~5 .lut_mask = 16'hDDA0;
defparam \Mux48~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N29
dffeas \reg_file[22][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][15] .is_wysiwyg = "true";
defparam \reg_file[22][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N21
dffeas \reg_file[18][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][15] .is_wysiwyg = "true";
defparam \reg_file[18][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N20
cycloneive_lcell_comb \Mux48~2 (
// Equation(s):
// \Mux48~2_combout  = (\prif.imemload_id [18] & ((\reg_file[22][15]~q ) # ((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (((\reg_file[18][15]~q  & !\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[22][15]~q ),
	.datac(\reg_file[18][15]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux48~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~2 .lut_mask = 16'hAAD8;
defparam \Mux48~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N19
dffeas \reg_file[30][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][15] .is_wysiwyg = "true";
defparam \reg_file[30][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N3
dffeas \reg_file[26][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][15] .is_wysiwyg = "true";
defparam \reg_file[26][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N18
cycloneive_lcell_comb \Mux48~3 (
// Equation(s):
// \Mux48~3_combout  = (\prif.imemload_id [19] & ((\Mux48~2_combout  & (\reg_file[30][15]~q )) # (!\Mux48~2_combout  & ((\reg_file[26][15]~q ))))) # (!\prif.imemload_id [19] & (\Mux48~2_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux48~2_combout ),
	.datac(\reg_file[30][15]~q ),
	.datad(\reg_file[26][15]~q ),
	.cin(gnd),
	.combout(\Mux48~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~3 .lut_mask = 16'hE6C4;
defparam \Mux48~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N10
cycloneive_lcell_comb \Mux48~6 (
// Equation(s):
// \Mux48~6_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16]) # (\Mux48~3_combout )))) # (!\prif.imemload_id [17] & (\Mux48~5_combout  & (!\prif.imemload_id [16])))

	.dataa(prifimemload_id_17),
	.datab(\Mux48~5_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux48~3_combout ),
	.cin(gnd),
	.combout(\Mux48~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~6 .lut_mask = 16'hAEA4;
defparam \Mux48~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N20
cycloneive_lcell_comb \reg_file[2][15]~feeder (
// Equation(s):
// \reg_file[2][15]~feeder_combout  = \reg_file_nxt[31][15]~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][15]~73_combout ),
	.cin(gnd),
	.combout(\reg_file[2][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][15]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[2][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y27_N21
dffeas \reg_file[2][15] (
	.clk(!CLK),
	.d(\reg_file[2][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][15] .is_wysiwyg = "true";
defparam \reg_file[2][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N30
cycloneive_lcell_comb \reg_file[3][15]~feeder (
// Equation(s):
// \reg_file[3][15]~feeder_combout  = \reg_file_nxt[31][15]~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][15]~73_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[3][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[3][15]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[3][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y27_N31
dffeas \reg_file[3][15] (
	.clk(!CLK),
	.d(\reg_file[3][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][15] .is_wysiwyg = "true";
defparam \reg_file[3][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N17
dffeas \reg_file[1][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][15] .is_wysiwyg = "true";
defparam \reg_file[1][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N26
cycloneive_lcell_comb \Mux48~14 (
// Equation(s):
// \Mux48~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][15]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][15]~q )))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[3][15]~q ),
	.datad(\reg_file[1][15]~q ),
	.cin(gnd),
	.combout(\Mux48~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~14 .lut_mask = 16'hC480;
defparam \Mux48~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N14
cycloneive_lcell_comb \Mux48~15 (
// Equation(s):
// \Mux48~15_combout  = (\Mux48~14_combout ) # ((!\prif.imemload_id [16] & (\reg_file[2][15]~q  & \prif.imemload_id [17])))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[2][15]~q ),
	.datac(prifimemload_id_17),
	.datad(\Mux48~14_combout ),
	.cin(gnd),
	.combout(\Mux48~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~15 .lut_mask = 16'hFF40;
defparam \Mux48~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N15
dffeas \reg_file[9][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][15] .is_wysiwyg = "true";
defparam \reg_file[9][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N29
dffeas \reg_file[11][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][15] .is_wysiwyg = "true";
defparam \reg_file[11][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N17
dffeas \reg_file[10][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][15] .is_wysiwyg = "true";
defparam \reg_file[10][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N15
dffeas \reg_file[8][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][15] .is_wysiwyg = "true";
defparam \reg_file[8][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N14
cycloneive_lcell_comb \Mux48~12 (
// Equation(s):
// \Mux48~12_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[10][15]~q )) # (!\prif.imemload_id [17] & ((\reg_file[8][15]~q )))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[10][15]~q ),
	.datac(\reg_file[8][15]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux48~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~12 .lut_mask = 16'hEE50;
defparam \Mux48~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N28
cycloneive_lcell_comb \Mux48~13 (
// Equation(s):
// \Mux48~13_combout  = (\prif.imemload_id [16] & ((\Mux48~12_combout  & ((\reg_file[11][15]~q ))) # (!\Mux48~12_combout  & (\reg_file[9][15]~q )))) # (!\prif.imemload_id [16] & (((\Mux48~12_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[9][15]~q ),
	.datac(\reg_file[11][15]~q ),
	.datad(\Mux48~12_combout ),
	.cin(gnd),
	.combout(\Mux48~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~13 .lut_mask = 16'hF588;
defparam \Mux48~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N6
cycloneive_lcell_comb \Mux48~16 (
// Equation(s):
// \Mux48~16_combout  = (\prif.imemload_id [19] & (((\Mux48~13_combout ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\Mux48~15_combout  & ((!\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\Mux48~15_combout ),
	.datac(\Mux48~13_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux48~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~16 .lut_mask = 16'hAAE4;
defparam \Mux48~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N6
cycloneive_lcell_comb \reg_file[6][15]~feeder (
// Equation(s):
// \reg_file[6][15]~feeder_combout  = \reg_file_nxt[31][15]~73_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][15]~73_combout ),
	.cin(gnd),
	.combout(\reg_file[6][15]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][15]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[6][15]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N7
dffeas \reg_file[6][15] (
	.clk(!CLK),
	.d(\reg_file[6][15]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][15] .is_wysiwyg = "true";
defparam \reg_file[6][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N31
dffeas \reg_file[5][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][15] .is_wysiwyg = "true";
defparam \reg_file[5][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N25
dffeas \reg_file[4][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][15] .is_wysiwyg = "true";
defparam \reg_file[4][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N30
cycloneive_lcell_comb \Mux48~10 (
// Equation(s):
// \Mux48~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][15]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][15]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][15]~q ),
	.datad(\reg_file[4][15]~q ),
	.cin(gnd),
	.combout(\Mux48~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~10 .lut_mask = 16'hB9A8;
defparam \Mux48~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N27
dffeas \reg_file[7][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][15] .is_wysiwyg = "true";
defparam \reg_file[7][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N28
cycloneive_lcell_comb \Mux48~11 (
// Equation(s):
// \Mux48~11_combout  = (\Mux48~10_combout  & (((\reg_file[7][15]~q ) # (!\prif.imemload_id [17])))) # (!\Mux48~10_combout  & (\reg_file[6][15]~q  & (\prif.imemload_id [17])))

	.dataa(\reg_file[6][15]~q ),
	.datab(\Mux48~10_combout ),
	.datac(prifimemload_id_17),
	.datad(\reg_file[7][15]~q ),
	.cin(gnd),
	.combout(\Mux48~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~11 .lut_mask = 16'hEC2C;
defparam \Mux48~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y26_N11
dffeas \reg_file[12][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][15] .is_wysiwyg = "true";
defparam \reg_file[12][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N13
dffeas \reg_file[13][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][15] .is_wysiwyg = "true";
defparam \reg_file[13][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N10
cycloneive_lcell_comb \Mux48~17 (
// Equation(s):
// \Mux48~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][15]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][15]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][15]~q ),
	.datad(\reg_file[13][15]~q ),
	.cin(gnd),
	.combout(\Mux48~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~17 .lut_mask = 16'hDC98;
defparam \Mux48~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y26_N25
dffeas \reg_file[14][15] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][15]~73_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][15] .is_wysiwyg = "true";
defparam \reg_file[14][15] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N27
dffeas \reg_file[15][15] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][15]~73_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][15]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][15] .is_wysiwyg = "true";
defparam \reg_file[15][15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N24
cycloneive_lcell_comb \Mux48~18 (
// Equation(s):
// \Mux48~18_combout  = (\prif.imemload_id [17] & ((\Mux48~17_combout  & ((\reg_file[15][15]~q ))) # (!\Mux48~17_combout  & (\reg_file[14][15]~q )))) # (!\prif.imemload_id [17] & (\Mux48~17_combout ))

	.dataa(prifimemload_id_17),
	.datab(\Mux48~17_combout ),
	.datac(\reg_file[14][15]~q ),
	.datad(\reg_file[15][15]~q ),
	.cin(gnd),
	.combout(\Mux48~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux48~18 .lut_mask = 16'hEC64;
defparam \Mux48~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N8
cycloneive_lcell_comb \reg_file_nxt[31][14]~74 (
// Equation(s):
// \reg_file_nxt[31][14]~74_combout  = (\Mux150~1_combout  & ((\prif.regwrite_wb [0]) # ((\prif.regwrite_wb [2]) # (!Equal8))))

	.dataa(prifregwrite_wb_0),
	.datab(prifregwrite_wb_2),
	.datac(Equal8),
	.datad(Mux150),
	.cin(gnd),
	.combout(\reg_file_nxt[31][14]~74_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][14]~74 .lut_mask = 16'hEF00;
defparam \reg_file_nxt[31][14]~74 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y30_N7
dffeas \reg_file[18][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][14] .is_wysiwyg = "true";
defparam \reg_file[18][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N22
cycloneive_lcell_comb \reg_file[26][14]~feeder (
// Equation(s):
// \reg_file[26][14]~feeder_combout  = \reg_file_nxt[31][14]~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][14]~74_combout ),
	.cin(gnd),
	.combout(\reg_file[26][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[26][14]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[26][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N23
dffeas \reg_file[26][14] (
	.clk(!CLK),
	.d(\reg_file[26][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][14] .is_wysiwyg = "true";
defparam \reg_file[26][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N6
cycloneive_lcell_comb \Mux49~2 (
// Equation(s):
// \Mux49~2_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[26][14]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & (\reg_file[18][14]~q )))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][14]~q ),
	.datad(\reg_file[26][14]~q ),
	.cin(gnd),
	.combout(\Mux49~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~2 .lut_mask = 16'hBA98;
defparam \Mux49~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N17
dffeas \reg_file[22][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][14] .is_wysiwyg = "true";
defparam \reg_file[22][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N20
cycloneive_lcell_comb \Mux49~3 (
// Equation(s):
// \Mux49~3_combout  = (\Mux49~2_combout  & ((\reg_file[30][14]~q ) # ((!\prif.imemload_id [18])))) # (!\Mux49~2_combout  & (((\prif.imemload_id [18] & \reg_file[22][14]~q ))))

	.dataa(\reg_file[30][14]~q ),
	.datab(\Mux49~2_combout ),
	.datac(prifimemload_id_18),
	.datad(\reg_file[22][14]~q ),
	.cin(gnd),
	.combout(\Mux49~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~3 .lut_mask = 16'hBC8C;
defparam \Mux49~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N9
dffeas \reg_file[28][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][14] .is_wysiwyg = "true";
defparam \reg_file[28][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N1
dffeas \reg_file[20][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][14] .is_wysiwyg = "true";
defparam \reg_file[20][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N7
dffeas \reg_file[16][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][14] .is_wysiwyg = "true";
defparam \reg_file[16][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y33_N11
dffeas \reg_file[24][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][14] .is_wysiwyg = "true";
defparam \reg_file[24][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N10
cycloneive_lcell_comb \Mux49~4 (
// Equation(s):
// \Mux49~4_combout  = (\prif.imemload_id [19] & (((\reg_file[24][14]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[16][14]~q  & ((!\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[16][14]~q ),
	.datac(\reg_file[24][14]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux49~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~4 .lut_mask = 16'hAAE4;
defparam \Mux49~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N0
cycloneive_lcell_comb \Mux49~5 (
// Equation(s):
// \Mux49~5_combout  = (\prif.imemload_id [18] & ((\Mux49~4_combout  & (\reg_file[28][14]~q )) # (!\Mux49~4_combout  & ((\reg_file[20][14]~q ))))) # (!\prif.imemload_id [18] & (((\Mux49~4_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[28][14]~q ),
	.datac(\reg_file[20][14]~q ),
	.datad(\Mux49~4_combout ),
	.cin(gnd),
	.combout(\Mux49~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~5 .lut_mask = 16'hDDA0;
defparam \Mux49~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N10
cycloneive_lcell_comb \Mux49~6 (
// Equation(s):
// \Mux49~6_combout  = (\prif.imemload_id [17] & ((\Mux49~3_combout ) # ((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (((\Mux49~5_combout  & !\prif.imemload_id [16]))))

	.dataa(prifimemload_id_17),
	.datab(\Mux49~3_combout ),
	.datac(\Mux49~5_combout ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux49~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~6 .lut_mask = 16'hAAD8;
defparam \Mux49~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y26_N7
dffeas \reg_file[23][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][14] .is_wysiwyg = "true";
defparam \reg_file[23][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N1
dffeas \reg_file[19][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][14] .is_wysiwyg = "true";
defparam \reg_file[19][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N6
cycloneive_lcell_comb \Mux49~7 (
// Equation(s):
// \Mux49~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][14]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][14]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][14]~q ),
	.datad(\reg_file[19][14]~q ),
	.cin(gnd),
	.combout(\Mux49~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~7 .lut_mask = 16'hB9A8;
defparam \Mux49~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N14
cycloneive_lcell_comb \reg_file[27][14]~feeder (
// Equation(s):
// \reg_file[27][14]~feeder_combout  = \reg_file_nxt[31][14]~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][14]~74_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[27][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[27][14]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[27][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N15
dffeas \reg_file[27][14] (
	.clk(!CLK),
	.d(\reg_file[27][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][14] .is_wysiwyg = "true";
defparam \reg_file[27][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N28
cycloneive_lcell_comb \reg_file[31][14]~feeder (
// Equation(s):
// \reg_file[31][14]~feeder_combout  = \reg_file_nxt[31][14]~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][14]~74_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[31][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][14]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[31][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y26_N29
dffeas \reg_file[31][14] (
	.clk(!CLK),
	.d(\reg_file[31][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][14] .is_wysiwyg = "true";
defparam \reg_file[31][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N0
cycloneive_lcell_comb \Mux49~8 (
// Equation(s):
// \Mux49~8_combout  = (\Mux49~7_combout  & (((\reg_file[31][14]~q ) # (!\prif.imemload_id [19])))) # (!\Mux49~7_combout  & (\reg_file[27][14]~q  & ((\prif.imemload_id [19]))))

	.dataa(\Mux49~7_combout ),
	.datab(\reg_file[27][14]~q ),
	.datac(\reg_file[31][14]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux49~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~8 .lut_mask = 16'hE4AA;
defparam \Mux49~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N8
cycloneive_lcell_comb \reg_file[25][14]~feeder (
// Equation(s):
// \reg_file[25][14]~feeder_combout  = \reg_file_nxt[31][14]~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][14]~74_combout ),
	.cin(gnd),
	.combout(\reg_file[25][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][14]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[25][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N9
dffeas \reg_file[25][14] (
	.clk(!CLK),
	.d(\reg_file[25][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][14] .is_wysiwyg = "true";
defparam \reg_file[25][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y28_N25
dffeas \reg_file[29][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][14] .is_wysiwyg = "true";
defparam \reg_file[29][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N29
dffeas \reg_file[17][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][14] .is_wysiwyg = "true";
defparam \reg_file[17][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N21
dffeas \reg_file[21][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][14] .is_wysiwyg = "true";
defparam \reg_file[21][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N20
cycloneive_lcell_comb \Mux49~0 (
// Equation(s):
// \Mux49~0_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[21][14]~q ))) # (!\prif.imemload_id [18] & (\reg_file[17][14]~q ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[17][14]~q ),
	.datac(\reg_file[21][14]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux49~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~0 .lut_mask = 16'hFA44;
defparam \Mux49~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N24
cycloneive_lcell_comb \Mux49~1 (
// Equation(s):
// \Mux49~1_combout  = (\prif.imemload_id [19] & ((\Mux49~0_combout  & ((\reg_file[29][14]~q ))) # (!\Mux49~0_combout  & (\reg_file[25][14]~q )))) # (!\prif.imemload_id [19] & (((\Mux49~0_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[25][14]~q ),
	.datac(\reg_file[29][14]~q ),
	.datad(\Mux49~0_combout ),
	.cin(gnd),
	.combout(\Mux49~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~1 .lut_mask = 16'hF588;
defparam \Mux49~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y26_N5
dffeas \reg_file[13][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][14] .is_wysiwyg = "true";
defparam \reg_file[13][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N27
dffeas \reg_file[12][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][14] .is_wysiwyg = "true";
defparam \reg_file[12][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N26
cycloneive_lcell_comb \Mux49~17 (
// Equation(s):
// \Mux49~17_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & (\reg_file[13][14]~q )) # (!\prif.imemload_id [16] & ((\reg_file[12][14]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[13][14]~q ),
	.datac(\reg_file[12][14]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux49~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~17 .lut_mask = 16'hEE50;
defparam \Mux49~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N9
dffeas \reg_file[15][14] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][14]~74_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][14] .is_wysiwyg = "true";
defparam \reg_file[15][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N14
cycloneive_lcell_comb \reg_file[14][14]~feeder (
// Equation(s):
// \reg_file[14][14]~feeder_combout  = \reg_file_nxt[31][14]~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][14]~74_combout ),
	.cin(gnd),
	.combout(\reg_file[14][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][14]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[14][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y26_N15
dffeas \reg_file[14][14] (
	.clk(!CLK),
	.d(\reg_file[14][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][14] .is_wysiwyg = "true";
defparam \reg_file[14][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N10
cycloneive_lcell_comb \Mux49~18 (
// Equation(s):
// \Mux49~18_combout  = (\Mux49~17_combout  & ((\reg_file[15][14]~q ) # ((!\prif.imemload_id [17])))) # (!\Mux49~17_combout  & (((\prif.imemload_id [17] & \reg_file[14][14]~q ))))

	.dataa(\Mux49~17_combout ),
	.datab(\reg_file[15][14]~q ),
	.datac(prifimemload_id_17),
	.datad(\reg_file[14][14]~q ),
	.cin(gnd),
	.combout(\Mux49~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~18 .lut_mask = 16'hDA8A;
defparam \Mux49~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N29
dffeas \reg_file[10][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][14] .is_wysiwyg = "true";
defparam \reg_file[10][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N28
cycloneive_lcell_comb \Mux49~10 (
// Equation(s):
// \Mux49~10_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][14]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][14]~q ))))

	.dataa(\reg_file[8][14]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[10][14]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux49~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~10 .lut_mask = 16'hFC22;
defparam \Mux49~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N26
cycloneive_lcell_comb \reg_file[9][14]~feeder (
// Equation(s):
// \reg_file[9][14]~feeder_combout  = \reg_file_nxt[31][14]~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][14]~74_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[9][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[9][14]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[9][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N27
dffeas \reg_file[9][14] (
	.clk(!CLK),
	.d(\reg_file[9][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][14] .is_wysiwyg = "true";
defparam \reg_file[9][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N13
dffeas \reg_file[11][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][14] .is_wysiwyg = "true";
defparam \reg_file[11][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N22
cycloneive_lcell_comb \Mux49~11 (
// Equation(s):
// \Mux49~11_combout  = (\prif.imemload_id [16] & ((\Mux49~10_combout  & ((\reg_file[11][14]~q ))) # (!\Mux49~10_combout  & (\reg_file[9][14]~q )))) # (!\prif.imemload_id [16] & (\Mux49~10_combout ))

	.dataa(prifimemload_id_16),
	.datab(\Mux49~10_combout ),
	.datac(\reg_file[9][14]~q ),
	.datad(\reg_file[11][14]~q ),
	.cin(gnd),
	.combout(\Mux49~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~11 .lut_mask = 16'hEC64;
defparam \Mux49~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N2
cycloneive_lcell_comb \reg_file[6][14]~feeder (
// Equation(s):
// \reg_file[6][14]~feeder_combout  = \reg_file_nxt[31][14]~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][14]~74_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][14]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y26_N3
dffeas \reg_file[6][14] (
	.clk(!CLK),
	.d(\reg_file[6][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][14] .is_wysiwyg = "true";
defparam \reg_file[6][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y32_N31
dffeas \reg_file[7][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][14] .is_wysiwyg = "true";
defparam \reg_file[7][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N27
dffeas \reg_file[4][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][14] .is_wysiwyg = "true";
defparam \reg_file[4][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N17
dffeas \reg_file[5][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][14] .is_wysiwyg = "true";
defparam \reg_file[5][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N26
cycloneive_lcell_comb \Mux49~12 (
// Equation(s):
// \Mux49~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][14]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][14]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][14]~q ),
	.datad(\reg_file[5][14]~q ),
	.cin(gnd),
	.combout(\Mux49~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~12 .lut_mask = 16'hBA98;
defparam \Mux49~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N30
cycloneive_lcell_comb \Mux49~13 (
// Equation(s):
// \Mux49~13_combout  = (\prif.imemload_id [17] & ((\Mux49~12_combout  & ((\reg_file[7][14]~q ))) # (!\Mux49~12_combout  & (\reg_file[6][14]~q )))) # (!\prif.imemload_id [17] & (((\Mux49~12_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][14]~q ),
	.datac(\reg_file[7][14]~q ),
	.datad(\Mux49~12_combout ),
	.cin(gnd),
	.combout(\Mux49~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~13 .lut_mask = 16'hF588;
defparam \Mux49~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N25
dffeas \reg_file[2][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][14] .is_wysiwyg = "true";
defparam \reg_file[2][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N7
dffeas \reg_file[1][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][14] .is_wysiwyg = "true";
defparam \reg_file[1][14] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y27_N21
dffeas \reg_file[3][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][14] .is_wysiwyg = "true";
defparam \reg_file[3][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N6
cycloneive_lcell_comb \Mux49~14 (
// Equation(s):
// \Mux49~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][14]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][14]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][14]~q ),
	.datad(\reg_file[3][14]~q ),
	.cin(gnd),
	.combout(\Mux49~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~14 .lut_mask = 16'hC840;
defparam \Mux49~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N24
cycloneive_lcell_comb \Mux49~15 (
// Equation(s):
// \Mux49~15_combout  = (\Mux49~14_combout ) # ((\prif.imemload_id [17] & (!\prif.imemload_id [16] & \reg_file[2][14]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[2][14]~q ),
	.datad(\Mux49~14_combout ),
	.cin(gnd),
	.combout(\Mux49~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~15 .lut_mask = 16'hFF20;
defparam \Mux49~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N22
cycloneive_lcell_comb \Mux49~16 (
// Equation(s):
// \Mux49~16_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\Mux49~13_combout )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\Mux49~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux49~13_combout ),
	.datad(\Mux49~15_combout ),
	.cin(gnd),
	.combout(\Mux49~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux49~16 .lut_mask = 16'hB9A8;
defparam \Mux49~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N16
cycloneive_lcell_comb \reg_file_nxt[31][13]~75 (
// Equation(s):
// \reg_file_nxt[31][13]~75_combout  = (\Mux151~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Mux151),
	.datac(prifregwrite_wb_0),
	.datad(Equal8),
	.cin(gnd),
	.combout(\reg_file_nxt[31][13]~75_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][13]~75 .lut_mask = 16'hC8CC;
defparam \reg_file_nxt[31][13]~75 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N15
dffeas \reg_file[30][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][13] .is_wysiwyg = "true";
defparam \reg_file[30][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N16
cycloneive_lcell_comb \reg_file[22][13]~feeder (
// Equation(s):
// \reg_file[22][13]~feeder_combout  = \reg_file_nxt[31][13]~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][13]~75_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[22][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][13]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[22][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N17
dffeas \reg_file[22][13] (
	.clk(!CLK),
	.d(\reg_file[22][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][13] .is_wysiwyg = "true";
defparam \reg_file[22][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N5
dffeas \reg_file[18][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][13] .is_wysiwyg = "true";
defparam \reg_file[18][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N4
cycloneive_lcell_comb \Mux50~2 (
// Equation(s):
// \Mux50~2_combout  = (\prif.imemload_id [18] & ((\reg_file[22][13]~q ) # ((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (((\reg_file[18][13]~q  & !\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[22][13]~q ),
	.datac(\reg_file[18][13]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux50~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~2 .lut_mask = 16'hAAD8;
defparam \Mux50~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N8
cycloneive_lcell_comb \Mux50~3 (
// Equation(s):
// \Mux50~3_combout  = (\prif.imemload_id [19] & ((\Mux50~2_combout  & ((\reg_file[30][13]~q ))) # (!\Mux50~2_combout  & (\reg_file[26][13]~q )))) # (!\prif.imemload_id [19] & (((\Mux50~2_combout ))))

	.dataa(\reg_file[26][13]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[30][13]~q ),
	.datad(\Mux50~2_combout ),
	.cin(gnd),
	.combout(\Mux50~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~3 .lut_mask = 16'hF388;
defparam \Mux50~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N23
dffeas \reg_file[24][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][13] .is_wysiwyg = "true";
defparam \reg_file[24][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N29
dffeas \reg_file[20][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][13] .is_wysiwyg = "true";
defparam \reg_file[20][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N28
cycloneive_lcell_comb \Mux50~4 (
// Equation(s):
// \Mux50~4_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[20][13]~q ))) # (!\prif.imemload_id [18] & (\reg_file[16][13]~q ))))

	.dataa(\reg_file[16][13]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[20][13]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux50~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~4 .lut_mask = 16'hFC22;
defparam \Mux50~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N22
cycloneive_lcell_comb \Mux50~5 (
// Equation(s):
// \Mux50~5_combout  = (\prif.imemload_id [19] & ((\Mux50~4_combout  & (\reg_file[28][13]~q )) # (!\Mux50~4_combout  & ((\reg_file[24][13]~q ))))) # (!\prif.imemload_id [19] & (((\Mux50~4_combout ))))

	.dataa(\reg_file[28][13]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[24][13]~q ),
	.datad(\Mux50~4_combout ),
	.cin(gnd),
	.combout(\Mux50~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~5 .lut_mask = 16'hBBC0;
defparam \Mux50~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N6
cycloneive_lcell_comb \Mux50~6 (
// Equation(s):
// \Mux50~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux50~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & ((\Mux50~5_combout ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux50~3_combout ),
	.datad(\Mux50~5_combout ),
	.cin(gnd),
	.combout(\Mux50~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~6 .lut_mask = 16'hB9A8;
defparam \Mux50~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y26_N19
dffeas \reg_file[25][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][13] .is_wysiwyg = "true";
defparam \reg_file[25][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N18
cycloneive_lcell_comb \Mux50~0 (
// Equation(s):
// \Mux50~0_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[25][13]~q ))) # (!\prif.imemload_id [19] & (\reg_file[17][13]~q ))))

	.dataa(\reg_file[17][13]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[25][13]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux50~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~0 .lut_mask = 16'hFC22;
defparam \Mux50~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y26_N21
dffeas \reg_file[21][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][13] .is_wysiwyg = "true";
defparam \reg_file[21][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N20
cycloneive_lcell_comb \reg_file[29][13]~feeder (
// Equation(s):
// \reg_file[29][13]~feeder_combout  = \reg_file_nxt[31][13]~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][13]~75_combout ),
	.cin(gnd),
	.combout(\reg_file[29][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][13]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N21
dffeas \reg_file[29][13] (
	.clk(!CLK),
	.d(\reg_file[29][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][13] .is_wysiwyg = "true";
defparam \reg_file[29][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N20
cycloneive_lcell_comb \Mux50~1 (
// Equation(s):
// \Mux50~1_combout  = (\prif.imemload_id [18] & ((\Mux50~0_combout  & ((\reg_file[29][13]~q ))) # (!\Mux50~0_combout  & (\reg_file[21][13]~q )))) # (!\prif.imemload_id [18] & (\Mux50~0_combout ))

	.dataa(prifimemload_id_18),
	.datab(\Mux50~0_combout ),
	.datac(\reg_file[21][13]~q ),
	.datad(\reg_file[29][13]~q ),
	.cin(gnd),
	.combout(\Mux50~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~1 .lut_mask = 16'hEC64;
defparam \Mux50~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y26_N21
dffeas \reg_file[31][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][13] .is_wysiwyg = "true";
defparam \reg_file[31][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N3
dffeas \reg_file[23][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][13] .is_wysiwyg = "true";
defparam \reg_file[23][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y26_N7
dffeas \reg_file[27][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][13] .is_wysiwyg = "true";
defparam \reg_file[27][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N25
dffeas \reg_file[19][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][13] .is_wysiwyg = "true";
defparam \reg_file[19][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N6
cycloneive_lcell_comb \Mux50~7 (
// Equation(s):
// \Mux50~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][13]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][13]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][13]~q ),
	.datad(\reg_file[19][13]~q ),
	.cin(gnd),
	.combout(\Mux50~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~7 .lut_mask = 16'hD9C8;
defparam \Mux50~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N2
cycloneive_lcell_comb \Mux50~8 (
// Equation(s):
// \Mux50~8_combout  = (\prif.imemload_id [18] & ((\Mux50~7_combout  & (\reg_file[31][13]~q )) # (!\Mux50~7_combout  & ((\reg_file[23][13]~q ))))) # (!\prif.imemload_id [18] & (((\Mux50~7_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[31][13]~q ),
	.datac(\reg_file[23][13]~q ),
	.datad(\Mux50~7_combout ),
	.cin(gnd),
	.combout(\Mux50~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~8 .lut_mask = 16'hDDA0;
defparam \Mux50~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N8
cycloneive_lcell_comb \reg_file[6][13]~feeder (
// Equation(s):
// \reg_file[6][13]~feeder_combout  = \reg_file_nxt[31][13]~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][13]~75_combout ),
	.cin(gnd),
	.combout(\reg_file[6][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][13]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[6][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y26_N9
dffeas \reg_file[6][13] (
	.clk(!CLK),
	.d(\reg_file[6][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][13] .is_wysiwyg = "true";
defparam \reg_file[6][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N19
dffeas \reg_file[7][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][13] .is_wysiwyg = "true";
defparam \reg_file[7][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N18
cycloneive_lcell_comb \reg_file[5][13]~feeder (
// Equation(s):
// \reg_file[5][13]~feeder_combout  = \reg_file_nxt[31][13]~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][13]~75_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[5][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[5][13]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[5][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N19
dffeas \reg_file[5][13] (
	.clk(!CLK),
	.d(\reg_file[5][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][13] .is_wysiwyg = "true";
defparam \reg_file[5][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N9
dffeas \reg_file[4][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][13] .is_wysiwyg = "true";
defparam \reg_file[4][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N4
cycloneive_lcell_comb \Mux50~10 (
// Equation(s):
// \Mux50~10_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & (\reg_file[5][13]~q )) # (!\prif.imemload_id [16] & ((\reg_file[4][13]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[5][13]~q ),
	.datac(\reg_file[4][13]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux50~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~10 .lut_mask = 16'hEE50;
defparam \Mux50~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N14
cycloneive_lcell_comb \Mux50~11 (
// Equation(s):
// \Mux50~11_combout  = (\prif.imemload_id [17] & ((\Mux50~10_combout  & ((\reg_file[7][13]~q ))) # (!\Mux50~10_combout  & (\reg_file[6][13]~q )))) # (!\prif.imemload_id [17] & (((\Mux50~10_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][13]~q ),
	.datac(\reg_file[7][13]~q ),
	.datad(\Mux50~10_combout ),
	.cin(gnd),
	.combout(\Mux50~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~11 .lut_mask = 16'hF588;
defparam \Mux50~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y26_N29
dffeas \reg_file[13][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][13] .is_wysiwyg = "true";
defparam \reg_file[13][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N28
cycloneive_lcell_comb \Mux50~17 (
// Equation(s):
// \Mux50~17_combout  = (\prif.imemload_id [16] & (((\reg_file[13][13]~q ) # (\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & (\reg_file[12][13]~q  & ((!\prif.imemload_id [17]))))

	.dataa(\reg_file[12][13]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[13][13]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux50~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~17 .lut_mask = 16'hCCE2;
defparam \Mux50~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N17
dffeas \reg_file[15][13] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][13]~75_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][13] .is_wysiwyg = "true";
defparam \reg_file[15][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y29_N1
dffeas \reg_file[14][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][13] .is_wysiwyg = "true";
defparam \reg_file[14][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N0
cycloneive_lcell_comb \Mux50~18 (
// Equation(s):
// \Mux50~18_combout  = (\Mux50~17_combout  & ((\reg_file[15][13]~q ) # ((!\prif.imemload_id [17])))) # (!\Mux50~17_combout  & (((\reg_file[14][13]~q  & \prif.imemload_id [17]))))

	.dataa(\Mux50~17_combout ),
	.datab(\reg_file[15][13]~q ),
	.datac(\reg_file[14][13]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux50~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~18 .lut_mask = 16'hD8AA;
defparam \Mux50~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N15
dffeas \reg_file[2][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][13] .is_wysiwyg = "true";
defparam \reg_file[2][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N5
dffeas \reg_file[3][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][13] .is_wysiwyg = "true";
defparam \reg_file[3][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N23
dffeas \reg_file[1][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][13] .is_wysiwyg = "true";
defparam \reg_file[1][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N22
cycloneive_lcell_comb \Mux50~14 (
// Equation(s):
// \Mux50~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][13]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][13]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[3][13]~q ),
	.datac(\reg_file[1][13]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux50~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~14 .lut_mask = 16'hD800;
defparam \Mux50~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N14
cycloneive_lcell_comb \Mux50~15 (
// Equation(s):
// \Mux50~15_combout  = (\Mux50~14_combout ) # ((\prif.imemload_id [17] & (!\prif.imemload_id [16] & \reg_file[2][13]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[2][13]~q ),
	.datad(\Mux50~14_combout ),
	.cin(gnd),
	.combout(\Mux50~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~15 .lut_mask = 16'hFF20;
defparam \Mux50~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N19
dffeas \reg_file[11][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][13] .is_wysiwyg = "true";
defparam \reg_file[11][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N21
dffeas \reg_file[9][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][13] .is_wysiwyg = "true";
defparam \reg_file[9][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N18
cycloneive_lcell_comb \Mux50~13 (
// Equation(s):
// \Mux50~13_combout  = (\Mux50~12_combout  & (((\reg_file[11][13]~q )) # (!\prif.imemload_id [16]))) # (!\Mux50~12_combout  & (\prif.imemload_id [16] & ((\reg_file[9][13]~q ))))

	.dataa(\Mux50~12_combout ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[11][13]~q ),
	.datad(\reg_file[9][13]~q ),
	.cin(gnd),
	.combout(\Mux50~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~13 .lut_mask = 16'hE6A2;
defparam \Mux50~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N16
cycloneive_lcell_comb \Mux50~16 (
// Equation(s):
// \Mux50~16_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\Mux50~13_combout ))) # (!\prif.imemload_id [19] & (\Mux50~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux50~15_combout ),
	.datad(\Mux50~13_combout ),
	.cin(gnd),
	.combout(\Mux50~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux50~16 .lut_mask = 16'hDC98;
defparam \Mux50~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N22
cycloneive_lcell_comb \reg_file_nxt[31][12]~76 (
// Equation(s):
// \reg_file_nxt[31][12]~76_combout  = (\Mux152~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Equal8),
	.datac(prifregwrite_wb_0),
	.datad(Mux152),
	.cin(gnd),
	.combout(\reg_file_nxt[31][12]~76_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][12]~76 .lut_mask = 16'hFB00;
defparam \reg_file_nxt[31][12]~76 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N12
cycloneive_lcell_comb \reg_file[27][12]~feeder (
// Equation(s):
// \reg_file[27][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[27][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[27][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[27][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N13
dffeas \reg_file[27][12] (
	.clk(!CLK),
	.d(\reg_file[27][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][12] .is_wysiwyg = "true";
defparam \reg_file[27][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N5
dffeas \reg_file[19][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][12] .is_wysiwyg = "true";
defparam \reg_file[19][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N11
dffeas \reg_file[23][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][12] .is_wysiwyg = "true";
defparam \reg_file[23][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N10
cycloneive_lcell_comb \Mux51~7 (
// Equation(s):
// \Mux51~7_combout  = (\prif.imemload_id [18] & (((\reg_file[23][12]~q ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\reg_file[19][12]~q  & ((!\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[19][12]~q ),
	.datac(\reg_file[23][12]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux51~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~7 .lut_mask = 16'hAAE4;
defparam \Mux51~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N4
cycloneive_lcell_comb \reg_file[31][12]~feeder (
// Equation(s):
// \reg_file[31][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[31][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[31][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y26_N5
dffeas \reg_file[31][12] (
	.clk(!CLK),
	.d(\reg_file[31][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][12] .is_wysiwyg = "true";
defparam \reg_file[31][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N26
cycloneive_lcell_comb \Mux51~8 (
// Equation(s):
// \Mux51~8_combout  = (\Mux51~7_combout  & (((\reg_file[31][12]~q ) # (!\prif.imemload_id [19])))) # (!\Mux51~7_combout  & (\reg_file[27][12]~q  & (\prif.imemload_id [19])))

	.dataa(\reg_file[27][12]~q ),
	.datab(\Mux51~7_combout ),
	.datac(prifimemload_id_19),
	.datad(\reg_file[31][12]~q ),
	.cin(gnd),
	.combout(\Mux51~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~8 .lut_mask = 16'hEC2C;
defparam \Mux51~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N9
dffeas \reg_file[30][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][12] .is_wysiwyg = "true";
defparam \reg_file[30][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N26
cycloneive_lcell_comb \reg_file[22][12]~feeder (
// Equation(s):
// \reg_file[22][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][12]~76_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[22][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][12]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[22][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N27
dffeas \reg_file[22][12] (
	.clk(!CLK),
	.d(\reg_file[22][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][12] .is_wysiwyg = "true";
defparam \reg_file[22][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N21
dffeas \reg_file[18][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][12] .is_wysiwyg = "true";
defparam \reg_file[18][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N10
cycloneive_lcell_comb \reg_file[26][12]~feeder (
// Equation(s):
// \reg_file[26][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[26][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[26][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[26][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N11
dffeas \reg_file[26][12] (
	.clk(!CLK),
	.d(\reg_file[26][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][12] .is_wysiwyg = "true";
defparam \reg_file[26][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N20
cycloneive_lcell_comb \Mux51~2 (
// Equation(s):
// \Mux51~2_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[26][12]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & (\reg_file[18][12]~q )))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][12]~q ),
	.datad(\reg_file[26][12]~q ),
	.cin(gnd),
	.combout(\Mux51~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~2 .lut_mask = 16'hBA98;
defparam \Mux51~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N0
cycloneive_lcell_comb \Mux51~3 (
// Equation(s):
// \Mux51~3_combout  = (\prif.imemload_id [18] & ((\Mux51~2_combout  & (\reg_file[30][12]~q )) # (!\Mux51~2_combout  & ((\reg_file[22][12]~q ))))) # (!\prif.imemload_id [18] & (((\Mux51~2_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[30][12]~q ),
	.datac(\reg_file[22][12]~q ),
	.datad(\Mux51~2_combout ),
	.cin(gnd),
	.combout(\Mux51~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~3 .lut_mask = 16'hDDA0;
defparam \Mux51~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N18
cycloneive_lcell_comb \reg_file[28][12]~feeder (
// Equation(s):
// \reg_file[28][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][12]~76_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[28][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[28][12]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[28][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N19
dffeas \reg_file[28][12] (
	.clk(!CLK),
	.d(\reg_file[28][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][12] .is_wysiwyg = "true";
defparam \reg_file[28][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N19
dffeas \reg_file[20][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][12] .is_wysiwyg = "true";
defparam \reg_file[20][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N21
dffeas \reg_file[16][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][12] .is_wysiwyg = "true";
defparam \reg_file[16][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y33_N3
dffeas \reg_file[24][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][12] .is_wysiwyg = "true";
defparam \reg_file[24][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N4
cycloneive_lcell_comb \Mux51~4 (
// Equation(s):
// \Mux51~4_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[24][12]~q ))) # (!\prif.imemload_id [19] & (\reg_file[16][12]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[16][12]~q ),
	.datad(\reg_file[24][12]~q ),
	.cin(gnd),
	.combout(\Mux51~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~4 .lut_mask = 16'hDC98;
defparam \Mux51~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N18
cycloneive_lcell_comb \Mux51~5 (
// Equation(s):
// \Mux51~5_combout  = (\prif.imemload_id [18] & ((\Mux51~4_combout  & (\reg_file[28][12]~q )) # (!\Mux51~4_combout  & ((\reg_file[20][12]~q ))))) # (!\prif.imemload_id [18] & (((\Mux51~4_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[28][12]~q ),
	.datac(\reg_file[20][12]~q ),
	.datad(\Mux51~4_combout ),
	.cin(gnd),
	.combout(\Mux51~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~5 .lut_mask = 16'hDDA0;
defparam \Mux51~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N22
cycloneive_lcell_comb \Mux51~6 (
// Equation(s):
// \Mux51~6_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\Mux51~3_combout )) # (!\prif.imemload_id [17] & ((\Mux51~5_combout )))))

	.dataa(\Mux51~3_combout ),
	.datab(\Mux51~5_combout ),
	.datac(prifimemload_id_16),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux51~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~6 .lut_mask = 16'hFA0C;
defparam \Mux51~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N2
cycloneive_lcell_comb \reg_file[29][12]~feeder (
// Equation(s):
// \reg_file[29][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[29][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N3
dffeas \reg_file[29][12] (
	.clk(!CLK),
	.d(\reg_file[29][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][12] .is_wysiwyg = "true";
defparam \reg_file[29][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N14
cycloneive_lcell_comb \reg_file[25][12]~feeder (
// Equation(s):
// \reg_file[25][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[25][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[25][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y28_N15
dffeas \reg_file[25][12] (
	.clk(!CLK),
	.d(\reg_file[25][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][12] .is_wysiwyg = "true";
defparam \reg_file[25][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N2
cycloneive_lcell_comb \reg_file[21][12]~feeder (
// Equation(s):
// \reg_file[21][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[21][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[21][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N3
dffeas \reg_file[21][12] (
	.clk(!CLK),
	.d(\reg_file[21][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][12] .is_wysiwyg = "true";
defparam \reg_file[21][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N25
dffeas \reg_file[17][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][12] .is_wysiwyg = "true";
defparam \reg_file[17][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N28
cycloneive_lcell_comb \Mux51~0 (
// Equation(s):
// \Mux51~0_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[21][12]~q )) # (!\prif.imemload_id [18] & ((\reg_file[17][12]~q )))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[21][12]~q ),
	.datac(\reg_file[17][12]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux51~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~0 .lut_mask = 16'hEE50;
defparam \Mux51~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N0
cycloneive_lcell_comb \Mux51~1 (
// Equation(s):
// \Mux51~1_combout  = (\prif.imemload_id [19] & ((\Mux51~0_combout  & (\reg_file[29][12]~q )) # (!\Mux51~0_combout  & ((\reg_file[25][12]~q ))))) # (!\prif.imemload_id [19] & (((\Mux51~0_combout ))))

	.dataa(\reg_file[29][12]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[25][12]~q ),
	.datad(\Mux51~0_combout ),
	.cin(gnd),
	.combout(\Mux51~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~1 .lut_mask = 16'hBBC0;
defparam \Mux51~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N23
dffeas \reg_file[11][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][12] .is_wysiwyg = "true";
defparam \reg_file[11][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N15
dffeas \reg_file[8][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][12] .is_wysiwyg = "true";
defparam \reg_file[8][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N5
dffeas \reg_file[10][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][12] .is_wysiwyg = "true";
defparam \reg_file[10][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N4
cycloneive_lcell_comb \Mux51~10 (
// Equation(s):
// \Mux51~10_combout  = (\prif.imemload_id [17] & (((\reg_file[10][12]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][12]~q  & ((!\prif.imemload_id [16]))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[8][12]~q ),
	.datac(\reg_file[10][12]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux51~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~10 .lut_mask = 16'hAAE4;
defparam \Mux51~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N5
dffeas \reg_file[9][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][12] .is_wysiwyg = "true";
defparam \reg_file[9][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N4
cycloneive_lcell_comb \Mux51~11 (
// Equation(s):
// \Mux51~11_combout  = (\Mux51~10_combout  & ((\reg_file[11][12]~q ) # ((!\prif.imemload_id [16])))) # (!\Mux51~10_combout  & (((\reg_file[9][12]~q  & \prif.imemload_id [16]))))

	.dataa(\reg_file[11][12]~q ),
	.datab(\Mux51~10_combout ),
	.datac(\reg_file[9][12]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux51~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~11 .lut_mask = 16'hB8CC;
defparam \Mux51~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y25_N3
dffeas \reg_file[3][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][12] .is_wysiwyg = "true";
defparam \reg_file[3][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y25_N13
dffeas \reg_file[1][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][12] .is_wysiwyg = "true";
defparam \reg_file[1][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N12
cycloneive_lcell_comb \Mux51~14 (
// Equation(s):
// \Mux51~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][12]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][12]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[3][12]~q ),
	.datac(\reg_file[1][12]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux51~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~14 .lut_mask = 16'hD800;
defparam \Mux51~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N16
cycloneive_lcell_comb \reg_file[2][12]~feeder (
// Equation(s):
// \reg_file[2][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[2][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[2][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y29_N17
dffeas \reg_file[2][12] (
	.clk(!CLK),
	.d(\reg_file[2][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][12] .is_wysiwyg = "true";
defparam \reg_file[2][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N26
cycloneive_lcell_comb \Mux51~15 (
// Equation(s):
// \Mux51~15_combout  = (\Mux51~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][12]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\Mux51~14_combout ),
	.datad(\reg_file[2][12]~q ),
	.cin(gnd),
	.combout(\Mux51~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~15 .lut_mask = 16'hF4F0;
defparam \Mux51~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N23
dffeas \reg_file[4][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][12] .is_wysiwyg = "true";
defparam \reg_file[4][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N21
dffeas \reg_file[5][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][12] .is_wysiwyg = "true";
defparam \reg_file[5][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N22
cycloneive_lcell_comb \Mux51~12 (
// Equation(s):
// \Mux51~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][12]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][12]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][12]~q ),
	.datad(\reg_file[5][12]~q ),
	.cin(gnd),
	.combout(\Mux51~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~12 .lut_mask = 16'hBA98;
defparam \Mux51~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N24
cycloneive_lcell_comb \reg_file[7][12]~feeder (
// Equation(s):
// \reg_file[7][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[7][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[7][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[7][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y29_N25
dffeas \reg_file[7][12] (
	.clk(!CLK),
	.d(\reg_file[7][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][12] .is_wysiwyg = "true";
defparam \reg_file[7][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N10
cycloneive_lcell_comb \Mux51~13 (
// Equation(s):
// \Mux51~13_combout  = (\prif.imemload_id [17] & ((\Mux51~12_combout  & ((\reg_file[7][12]~q ))) # (!\Mux51~12_combout  & (\reg_file[6][12]~q )))) # (!\prif.imemload_id [17] & (((\Mux51~12_combout ))))

	.dataa(\reg_file[6][12]~q ),
	.datab(prifimemload_id_17),
	.datac(\Mux51~12_combout ),
	.datad(\reg_file[7][12]~q ),
	.cin(gnd),
	.combout(\Mux51~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~13 .lut_mask = 16'hF838;
defparam \Mux51~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N8
cycloneive_lcell_comb \Mux51~16 (
// Equation(s):
// \Mux51~16_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\Mux51~13_combout ))) # (!\prif.imemload_id [18] & (\Mux51~15_combout ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\Mux51~15_combout ),
	.datad(\Mux51~13_combout ),
	.cin(gnd),
	.combout(\Mux51~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~16 .lut_mask = 16'hDC98;
defparam \Mux51~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y26_N15
dffeas \reg_file[12][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][12] .is_wysiwyg = "true";
defparam \reg_file[12][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N1
dffeas \reg_file[13][12] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][12]~76_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][12] .is_wysiwyg = "true";
defparam \reg_file[13][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N14
cycloneive_lcell_comb \Mux51~17 (
// Equation(s):
// \Mux51~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][12]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][12]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][12]~q ),
	.datad(\reg_file[13][12]~q ),
	.cin(gnd),
	.combout(\Mux51~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~17 .lut_mask = 16'hDC98;
defparam \Mux51~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N22
cycloneive_lcell_comb \reg_file[14][12]~feeder (
// Equation(s):
// \reg_file[14][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[14][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[14][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N23
dffeas \reg_file[14][12] (
	.clk(!CLK),
	.d(\reg_file[14][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][12] .is_wysiwyg = "true";
defparam \reg_file[14][12] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N23
dffeas \reg_file[15][12] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][12]~76_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][12] .is_wysiwyg = "true";
defparam \reg_file[15][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N28
cycloneive_lcell_comb \Mux51~18 (
// Equation(s):
// \Mux51~18_combout  = (\prif.imemload_id [17] & ((\Mux51~17_combout  & ((\reg_file[15][12]~q ))) # (!\Mux51~17_combout  & (\reg_file[14][12]~q )))) # (!\prif.imemload_id [17] & (\Mux51~17_combout ))

	.dataa(prifimemload_id_17),
	.datab(\Mux51~17_combout ),
	.datac(\reg_file[14][12]~q ),
	.datad(\reg_file[15][12]~q ),
	.cin(gnd),
	.combout(\Mux51~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux51~18 .lut_mask = 16'hEC64;
defparam \Mux51~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N12
cycloneive_lcell_comb \reg_file_nxt[31][11]~77 (
// Equation(s):
// \reg_file_nxt[31][11]~77_combout  = (\Mux153~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Mux153),
	.datac(prifregwrite_wb_0),
	.datad(Equal8),
	.cin(gnd),
	.combout(\reg_file_nxt[31][11]~77_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][11]~77 .lut_mask = 16'hC8CC;
defparam \reg_file_nxt[31][11]~77 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N22
cycloneive_lcell_comb \reg_file[23][11]~feeder (
// Equation(s):
// \reg_file[23][11]~feeder_combout  = \reg_file_nxt[31][11]~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][11]~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[23][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][11]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[23][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y26_N23
dffeas \reg_file[23][11] (
	.clk(!CLK),
	.d(\reg_file[23][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][11] .is_wysiwyg = "true";
defparam \reg_file[23][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N17
dffeas \reg_file[31][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][11] .is_wysiwyg = "true";
defparam \reg_file[31][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y26_N11
dffeas \reg_file[27][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][11] .is_wysiwyg = "true";
defparam \reg_file[27][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N29
dffeas \reg_file[19][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][11] .is_wysiwyg = "true";
defparam \reg_file[19][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N10
cycloneive_lcell_comb \Mux52~7 (
// Equation(s):
// \Mux52~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][11]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][11]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][11]~q ),
	.datad(\reg_file[19][11]~q ),
	.cin(gnd),
	.combout(\Mux52~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~7 .lut_mask = 16'hD9C8;
defparam \Mux52~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N16
cycloneive_lcell_comb \Mux52~8 (
// Equation(s):
// \Mux52~8_combout  = (\prif.imemload_id [18] & ((\Mux52~7_combout  & ((\reg_file[31][11]~q ))) # (!\Mux52~7_combout  & (\reg_file[23][11]~q )))) # (!\prif.imemload_id [18] & (((\Mux52~7_combout ))))

	.dataa(\reg_file[23][11]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[31][11]~q ),
	.datad(\Mux52~7_combout ),
	.cin(gnd),
	.combout(\Mux52~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~8 .lut_mask = 16'hF388;
defparam \Mux52~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y26_N15
dffeas \reg_file[25][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][11] .is_wysiwyg = "true";
defparam \reg_file[25][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N14
cycloneive_lcell_comb \Mux52~0 (
// Equation(s):
// \Mux52~0_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[25][11]~q ))) # (!\prif.imemload_id [19] & (\reg_file[17][11]~q ))))

	.dataa(\reg_file[17][11]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[25][11]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux52~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~0 .lut_mask = 16'hFC22;
defparam \Mux52~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y26_N25
dffeas \reg_file[21][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][11] .is_wysiwyg = "true";
defparam \reg_file[21][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y29_N11
dffeas \reg_file[29][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][11] .is_wysiwyg = "true";
defparam \reg_file[29][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N24
cycloneive_lcell_comb \Mux52~1 (
// Equation(s):
// \Mux52~1_combout  = (\prif.imemload_id [18] & ((\Mux52~0_combout  & ((\reg_file[29][11]~q ))) # (!\Mux52~0_combout  & (\reg_file[21][11]~q )))) # (!\prif.imemload_id [18] & (\Mux52~0_combout ))

	.dataa(prifimemload_id_18),
	.datab(\Mux52~0_combout ),
	.datac(\reg_file[21][11]~q ),
	.datad(\reg_file[29][11]~q ),
	.cin(gnd),
	.combout(\Mux52~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~1 .lut_mask = 16'hEC64;
defparam \Mux52~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N9
dffeas \reg_file[28][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][11] .is_wysiwyg = "true";
defparam \reg_file[28][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N31
dffeas \reg_file[24][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][11] .is_wysiwyg = "true";
defparam \reg_file[24][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N15
dffeas \reg_file[16][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][11] .is_wysiwyg = "true";
defparam \reg_file[16][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N17
dffeas \reg_file[20][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][11] .is_wysiwyg = "true";
defparam \reg_file[20][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N16
cycloneive_lcell_comb \Mux52~4 (
// Equation(s):
// \Mux52~4_combout  = (\prif.imemload_id [18] & (((\reg_file[20][11]~q ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\reg_file[16][11]~q  & ((!\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[16][11]~q ),
	.datac(\reg_file[20][11]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux52~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~4 .lut_mask = 16'hAAE4;
defparam \Mux52~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N30
cycloneive_lcell_comb \Mux52~5 (
// Equation(s):
// \Mux52~5_combout  = (\prif.imemload_id [19] & ((\Mux52~4_combout  & (\reg_file[28][11]~q )) # (!\Mux52~4_combout  & ((\reg_file[24][11]~q ))))) # (!\prif.imemload_id [19] & (((\Mux52~4_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[28][11]~q ),
	.datac(\reg_file[24][11]~q ),
	.datad(\Mux52~4_combout ),
	.cin(gnd),
	.combout(\Mux52~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~5 .lut_mask = 16'hDDA0;
defparam \Mux52~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N31
dffeas \reg_file[26][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][11] .is_wysiwyg = "true";
defparam \reg_file[26][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N3
dffeas \reg_file[30][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][11] .is_wysiwyg = "true";
defparam \reg_file[30][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N29
dffeas \reg_file[18][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][11] .is_wysiwyg = "true";
defparam \reg_file[18][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N0
cycloneive_lcell_comb \reg_file[22][11]~feeder (
// Equation(s):
// \reg_file[22][11]~feeder_combout  = \reg_file_nxt[31][11]~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][11]~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[22][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][11]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[22][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N1
dffeas \reg_file[22][11] (
	.clk(!CLK),
	.d(\reg_file[22][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][11] .is_wysiwyg = "true";
defparam \reg_file[22][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N28
cycloneive_lcell_comb \Mux52~2 (
// Equation(s):
// \Mux52~2_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[22][11]~q ))) # (!\prif.imemload_id [18] & (\reg_file[18][11]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][11]~q ),
	.datad(\reg_file[22][11]~q ),
	.cin(gnd),
	.combout(\Mux52~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~2 .lut_mask = 16'hDC98;
defparam \Mux52~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N28
cycloneive_lcell_comb \Mux52~3 (
// Equation(s):
// \Mux52~3_combout  = (\prif.imemload_id [19] & ((\Mux52~2_combout  & ((\reg_file[30][11]~q ))) # (!\Mux52~2_combout  & (\reg_file[26][11]~q )))) # (!\prif.imemload_id [19] & (((\Mux52~2_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[26][11]~q ),
	.datac(\reg_file[30][11]~q ),
	.datad(\Mux52~2_combout ),
	.cin(gnd),
	.combout(\Mux52~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~3 .lut_mask = 16'hF588;
defparam \Mux52~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N6
cycloneive_lcell_comb \Mux52~6 (
// Equation(s):
// \Mux52~6_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\Mux52~3_combout ))) # (!\prif.imemload_id [17] & (\Mux52~5_combout ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\Mux52~5_combout ),
	.datad(\Mux52~3_combout ),
	.cin(gnd),
	.combout(\Mux52~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~6 .lut_mask = 16'hDC98;
defparam \Mux52~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N27
dffeas \reg_file[11][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][11] .is_wysiwyg = "true";
defparam \reg_file[11][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N25
dffeas \reg_file[9][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][11] .is_wysiwyg = "true";
defparam \reg_file[9][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N26
cycloneive_lcell_comb \Mux52~13 (
// Equation(s):
// \Mux52~13_combout  = (\Mux52~12_combout  & (((\reg_file[11][11]~q )) # (!\prif.imemload_id [16]))) # (!\Mux52~12_combout  & (\prif.imemload_id [16] & ((\reg_file[9][11]~q ))))

	.dataa(\Mux52~12_combout ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[11][11]~q ),
	.datad(\reg_file[9][11]~q ),
	.cin(gnd),
	.combout(\Mux52~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~13 .lut_mask = 16'hE6A2;
defparam \Mux52~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y29_N19
dffeas \reg_file[2][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][11] .is_wysiwyg = "true";
defparam \reg_file[2][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N29
dffeas \reg_file[3][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][11] .is_wysiwyg = "true";
defparam \reg_file[3][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N15
dffeas \reg_file[1][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][11] .is_wysiwyg = "true";
defparam \reg_file[1][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N28
cycloneive_lcell_comb \Mux52~14 (
// Equation(s):
// \Mux52~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][11]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][11]~q )))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[3][11]~q ),
	.datad(\reg_file[1][11]~q ),
	.cin(gnd),
	.combout(\Mux52~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~14 .lut_mask = 16'hC480;
defparam \Mux52~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N18
cycloneive_lcell_comb \Mux52~15 (
// Equation(s):
// \Mux52~15_combout  = (\Mux52~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][11]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[2][11]~q ),
	.datad(\Mux52~14_combout ),
	.cin(gnd),
	.combout(\Mux52~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~15 .lut_mask = 16'hFF40;
defparam \Mux52~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N20
cycloneive_lcell_comb \Mux52~16 (
// Equation(s):
// \Mux52~16_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\Mux52~13_combout )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & ((\Mux52~15_combout ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\Mux52~13_combout ),
	.datad(\Mux52~15_combout ),
	.cin(gnd),
	.combout(\Mux52~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~16 .lut_mask = 16'hB9A8;
defparam \Mux52~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N20
cycloneive_lcell_comb \reg_file[6][11]~feeder (
// Equation(s):
// \reg_file[6][11]~feeder_combout  = \reg_file_nxt[31][11]~77_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][11]~77_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][11]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][11]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][11]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y26_N21
dffeas \reg_file[6][11] (
	.clk(!CLK),
	.d(\reg_file[6][11]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][11] .is_wysiwyg = "true";
defparam \reg_file[6][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N29
dffeas \reg_file[4][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][11] .is_wysiwyg = "true";
defparam \reg_file[4][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N11
dffeas \reg_file[5][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][11] .is_wysiwyg = "true";
defparam \reg_file[5][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N10
cycloneive_lcell_comb \Mux52~10 (
// Equation(s):
// \Mux52~10_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[5][11]~q ))) # (!\prif.imemload_id [16] & (\reg_file[4][11]~q ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[4][11]~q ),
	.datac(\reg_file[5][11]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux52~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~10 .lut_mask = 16'hFA44;
defparam \Mux52~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N7
dffeas \reg_file[7][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][11] .is_wysiwyg = "true";
defparam \reg_file[7][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N6
cycloneive_lcell_comb \Mux52~11 (
// Equation(s):
// \Mux52~11_combout  = (\prif.imemload_id [17] & ((\Mux52~10_combout  & ((\reg_file[7][11]~q ))) # (!\Mux52~10_combout  & (\reg_file[6][11]~q )))) # (!\prif.imemload_id [17] & (((\Mux52~10_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][11]~q ),
	.datac(\Mux52~10_combout ),
	.datad(\reg_file[7][11]~q ),
	.cin(gnd),
	.combout(\Mux52~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~11 .lut_mask = 16'hF858;
defparam \Mux52~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N5
dffeas \reg_file[13][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][11] .is_wysiwyg = "true";
defparam \reg_file[13][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N19
dffeas \reg_file[12][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][11] .is_wysiwyg = "true";
defparam \reg_file[12][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N4
cycloneive_lcell_comb \Mux52~17 (
// Equation(s):
// \Mux52~17_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[13][11]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[12][11]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[13][11]~q ),
	.datad(\reg_file[12][11]~q ),
	.cin(gnd),
	.combout(\Mux52~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~17 .lut_mask = 16'hB9A8;
defparam \Mux52~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y26_N29
dffeas \reg_file[14][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][11] .is_wysiwyg = "true";
defparam \reg_file[14][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N13
dffeas \reg_file[15][11] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][11]~77_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][11] .is_wysiwyg = "true";
defparam \reg_file[15][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N28
cycloneive_lcell_comb \Mux52~18 (
// Equation(s):
// \Mux52~18_combout  = (\prif.imemload_id [17] & ((\Mux52~17_combout  & ((\reg_file[15][11]~q ))) # (!\Mux52~17_combout  & (\reg_file[14][11]~q )))) # (!\prif.imemload_id [17] & (\Mux52~17_combout ))

	.dataa(prifimemload_id_17),
	.datab(\Mux52~17_combout ),
	.datac(\reg_file[14][11]~q ),
	.datad(\reg_file[15][11]~q ),
	.cin(gnd),
	.combout(\Mux52~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux52~18 .lut_mask = 16'hEC64;
defparam \Mux52~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N2
cycloneive_lcell_comb \reg_file_nxt[31][10]~78 (
// Equation(s):
// \reg_file_nxt[31][10]~78_combout  = (\Mux154~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Mux154),
	.datac(prifregwrite_wb_0),
	.datad(Equal8),
	.cin(gnd),
	.combout(\reg_file_nxt[31][10]~78_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][10]~78 .lut_mask = 16'hC8CC;
defparam \reg_file_nxt[31][10]~78 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N21
dffeas \reg_file[29][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][10] .is_wysiwyg = "true";
defparam \reg_file[29][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y26_N1
dffeas \reg_file[25][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][10] .is_wysiwyg = "true";
defparam \reg_file[25][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N9
dffeas \reg_file[17][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][10] .is_wysiwyg = "true";
defparam \reg_file[17][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N10
cycloneive_lcell_comb \reg_file[21][10]~feeder (
// Equation(s):
// \reg_file[21][10]~feeder_combout  = \reg_file_nxt[31][10]~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][10]~78_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[21][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][10]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[21][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y26_N11
dffeas \reg_file[21][10] (
	.clk(!CLK),
	.d(\reg_file[21][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][10] .is_wysiwyg = "true";
defparam \reg_file[21][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N28
cycloneive_lcell_comb \Mux53~0 (
// Equation(s):
// \Mux53~0_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[21][10]~q ))) # (!\prif.imemload_id [18] & (\reg_file[17][10]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[17][10]~q ),
	.datad(\reg_file[21][10]~q ),
	.cin(gnd),
	.combout(\Mux53~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~0 .lut_mask = 16'hDC98;
defparam \Mux53~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N0
cycloneive_lcell_comb \Mux53~1 (
// Equation(s):
// \Mux53~1_combout  = (\prif.imemload_id [19] & ((\Mux53~0_combout  & (\reg_file[29][10]~q )) # (!\Mux53~0_combout  & ((\reg_file[25][10]~q ))))) # (!\prif.imemload_id [19] & (((\Mux53~0_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[29][10]~q ),
	.datac(\reg_file[25][10]~q ),
	.datad(\Mux53~0_combout ),
	.cin(gnd),
	.combout(\Mux53~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~1 .lut_mask = 16'hDDA0;
defparam \Mux53~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N25
dffeas \reg_file[18][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][10] .is_wysiwyg = "true";
defparam \reg_file[18][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N3
dffeas \reg_file[26][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][10] .is_wysiwyg = "true";
defparam \reg_file[26][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N24
cycloneive_lcell_comb \Mux53~2 (
// Equation(s):
// \Mux53~2_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[26][10]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & (\reg_file[18][10]~q )))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][10]~q ),
	.datad(\reg_file[26][10]~q ),
	.cin(gnd),
	.combout(\Mux53~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~2 .lut_mask = 16'hBA98;
defparam \Mux53~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N1
dffeas \reg_file[30][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][10] .is_wysiwyg = "true";
defparam \reg_file[30][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y30_N19
dffeas \reg_file[22][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][10] .is_wysiwyg = "true";
defparam \reg_file[22][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N0
cycloneive_lcell_comb \Mux53~3 (
// Equation(s):
// \Mux53~3_combout  = (\prif.imemload_id [18] & ((\Mux53~2_combout  & (\reg_file[30][10]~q )) # (!\Mux53~2_combout  & ((\reg_file[22][10]~q ))))) # (!\prif.imemload_id [18] & (\Mux53~2_combout ))

	.dataa(prifimemload_id_18),
	.datab(\Mux53~2_combout ),
	.datac(\reg_file[30][10]~q ),
	.datad(\reg_file[22][10]~q ),
	.cin(gnd),
	.combout(\Mux53~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~3 .lut_mask = 16'hE6C4;
defparam \Mux53~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N29
dffeas \reg_file[24][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][10] .is_wysiwyg = "true";
defparam \reg_file[24][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N5
dffeas \reg_file[16][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][10] .is_wysiwyg = "true";
defparam \reg_file[16][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N28
cycloneive_lcell_comb \Mux53~4 (
// Equation(s):
// \Mux53~4_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[24][10]~q )) # (!\prif.imemload_id [19] & ((\reg_file[16][10]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[24][10]~q ),
	.datad(\reg_file[16][10]~q ),
	.cin(gnd),
	.combout(\Mux53~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~4 .lut_mask = 16'hD9C8;
defparam \Mux53~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N11
dffeas \reg_file[20][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][10] .is_wysiwyg = "true";
defparam \reg_file[20][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N10
cycloneive_lcell_comb \Mux53~5 (
// Equation(s):
// \Mux53~5_combout  = (\Mux53~4_combout  & ((\reg_file[28][10]~q ) # ((!\prif.imemload_id [18])))) # (!\Mux53~4_combout  & (((\reg_file[20][10]~q  & \prif.imemload_id [18]))))

	.dataa(\reg_file[28][10]~q ),
	.datab(\Mux53~4_combout ),
	.datac(\reg_file[20][10]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux53~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~5 .lut_mask = 16'hB8CC;
defparam \Mux53~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N14
cycloneive_lcell_comb \Mux53~6 (
// Equation(s):
// \Mux53~6_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\Mux53~3_combout )) # (!\prif.imemload_id [17] & ((\Mux53~5_combout )))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\Mux53~3_combout ),
	.datad(\Mux53~5_combout ),
	.cin(gnd),
	.combout(\Mux53~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~6 .lut_mask = 16'hD9C8;
defparam \Mux53~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N18
cycloneive_lcell_comb \reg_file[27][10]~feeder (
// Equation(s):
// \reg_file[27][10]~feeder_combout  = \reg_file_nxt[31][10]~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][10]~78_combout ),
	.cin(gnd),
	.combout(\reg_file[27][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[27][10]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[27][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N19
dffeas \reg_file[27][10] (
	.clk(!CLK),
	.d(\reg_file[27][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][10] .is_wysiwyg = "true";
defparam \reg_file[27][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N27
dffeas \reg_file[31][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][10] .is_wysiwyg = "true";
defparam \reg_file[31][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N15
dffeas \reg_file[23][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][10] .is_wysiwyg = "true";
defparam \reg_file[23][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N21
dffeas \reg_file[19][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][10] .is_wysiwyg = "true";
defparam \reg_file[19][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N14
cycloneive_lcell_comb \Mux53~7 (
// Equation(s):
// \Mux53~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][10]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][10]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][10]~q ),
	.datad(\reg_file[19][10]~q ),
	.cin(gnd),
	.combout(\Mux53~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~7 .lut_mask = 16'hB9A8;
defparam \Mux53~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N26
cycloneive_lcell_comb \Mux53~8 (
// Equation(s):
// \Mux53~8_combout  = (\prif.imemload_id [19] & ((\Mux53~7_combout  & ((\reg_file[31][10]~q ))) # (!\Mux53~7_combout  & (\reg_file[27][10]~q )))) # (!\prif.imemload_id [19] & (((\Mux53~7_combout ))))

	.dataa(\reg_file[27][10]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[31][10]~q ),
	.datad(\Mux53~7_combout ),
	.cin(gnd),
	.combout(\Mux53~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~8 .lut_mask = 16'hF388;
defparam \Mux53~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N11
dffeas \reg_file[12][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][10] .is_wysiwyg = "true";
defparam \reg_file[12][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N17
dffeas \reg_file[13][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][10] .is_wysiwyg = "true";
defparam \reg_file[13][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N10
cycloneive_lcell_comb \Mux53~17 (
// Equation(s):
// \Mux53~17_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[13][10]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[12][10]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[12][10]~q ),
	.datad(\reg_file[13][10]~q ),
	.cin(gnd),
	.combout(\Mux53~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~17 .lut_mask = 16'hBA98;
defparam \Mux53~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N3
dffeas \reg_file[15][10] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][10]~78_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][10] .is_wysiwyg = "true";
defparam \reg_file[15][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N6
cycloneive_lcell_comb \reg_file[14][10]~feeder (
// Equation(s):
// \reg_file[14][10]~feeder_combout  = \reg_file_nxt[31][10]~78_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][10]~78_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[14][10]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][10]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[14][10]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N7
dffeas \reg_file[14][10] (
	.clk(!CLK),
	.d(\reg_file[14][10]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][10] .is_wysiwyg = "true";
defparam \reg_file[14][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N24
cycloneive_lcell_comb \Mux53~18 (
// Equation(s):
// \Mux53~18_combout  = (\Mux53~17_combout  & ((\reg_file[15][10]~q ) # ((!\prif.imemload_id [17])))) # (!\Mux53~17_combout  & (((\prif.imemload_id [17] & \reg_file[14][10]~q ))))

	.dataa(\Mux53~17_combout ),
	.datab(\reg_file[15][10]~q ),
	.datac(prifimemload_id_17),
	.datad(\reg_file[14][10]~q ),
	.cin(gnd),
	.combout(\Mux53~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~18 .lut_mask = 16'hDA8A;
defparam \Mux53~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N3
dffeas \reg_file[8][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][10] .is_wysiwyg = "true";
defparam \reg_file[8][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N13
dffeas \reg_file[10][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][10] .is_wysiwyg = "true";
defparam \reg_file[10][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N12
cycloneive_lcell_comb \Mux53~10 (
// Equation(s):
// \Mux53~10_combout  = (\prif.imemload_id [17] & (((\reg_file[10][10]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][10]~q  & ((!\prif.imemload_id [16]))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[8][10]~q ),
	.datac(\reg_file[10][10]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux53~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~10 .lut_mask = 16'hAAE4;
defparam \Mux53~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N29
dffeas \reg_file[9][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][10] .is_wysiwyg = "true";
defparam \reg_file[9][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N3
dffeas \reg_file[11][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][10] .is_wysiwyg = "true";
defparam \reg_file[11][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N28
cycloneive_lcell_comb \Mux53~11 (
// Equation(s):
// \Mux53~11_combout  = (\Mux53~10_combout  & (((\reg_file[11][10]~q )) # (!\prif.imemload_id [16]))) # (!\Mux53~10_combout  & (\prif.imemload_id [16] & (\reg_file[9][10]~q )))

	.dataa(\Mux53~10_combout ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[9][10]~q ),
	.datad(\reg_file[11][10]~q ),
	.cin(gnd),
	.combout(\Mux53~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~11 .lut_mask = 16'hEA62;
defparam \Mux53~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y29_N3
dffeas \reg_file[2][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][10] .is_wysiwyg = "true";
defparam \reg_file[2][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y25_N1
dffeas \reg_file[1][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][10] .is_wysiwyg = "true";
defparam \reg_file[1][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y25_N11
dffeas \reg_file[3][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][10] .is_wysiwyg = "true";
defparam \reg_file[3][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N10
cycloneive_lcell_comb \Mux53~14 (
// Equation(s):
// \Mux53~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][10]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][10]~q ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[1][10]~q ),
	.datac(\reg_file[3][10]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux53~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~14 .lut_mask = 16'hE400;
defparam \Mux53~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y29_N2
cycloneive_lcell_comb \Mux53~15 (
// Equation(s):
// \Mux53~15_combout  = (\Mux53~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][10]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[2][10]~q ),
	.datad(\Mux53~14_combout ),
	.cin(gnd),
	.combout(\Mux53~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~15 .lut_mask = 16'hFF40;
defparam \Mux53~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N25
dffeas \reg_file[6][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][10] .is_wysiwyg = "true";
defparam \reg_file[6][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N7
dffeas \reg_file[7][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][10] .is_wysiwyg = "true";
defparam \reg_file[7][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N5
dffeas \reg_file[5][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][10] .is_wysiwyg = "true";
defparam \reg_file[5][10] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N3
dffeas \reg_file[4][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][10] .is_wysiwyg = "true";
defparam \reg_file[4][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N4
cycloneive_lcell_comb \Mux53~12 (
// Equation(s):
// \Mux53~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][10]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][10]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][10]~q ),
	.datad(\reg_file[4][10]~q ),
	.cin(gnd),
	.combout(\Mux53~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~12 .lut_mask = 16'hB9A8;
defparam \Mux53~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N6
cycloneive_lcell_comb \Mux53~13 (
// Equation(s):
// \Mux53~13_combout  = (\prif.imemload_id [17] & ((\Mux53~12_combout  & ((\reg_file[7][10]~q ))) # (!\Mux53~12_combout  & (\reg_file[6][10]~q )))) # (!\prif.imemload_id [17] & (((\Mux53~12_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][10]~q ),
	.datac(\reg_file[7][10]~q ),
	.datad(\Mux53~12_combout ),
	.cin(gnd),
	.combout(\Mux53~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~13 .lut_mask = 16'hF588;
defparam \Mux53~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N16
cycloneive_lcell_comb \Mux53~16 (
// Equation(s):
// \Mux53~16_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\Mux53~13_combout ))) # (!\prif.imemload_id [18] & (\Mux53~15_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\Mux53~15_combout ),
	.datac(\Mux53~13_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux53~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux53~16 .lut_mask = 16'hFA44;
defparam \Mux53~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N10
cycloneive_lcell_comb \reg_file_nxt[31][9]~79 (
// Equation(s):
// \reg_file_nxt[31][9]~79_combout  = (\Mux155~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Equal8),
	.datac(prifregwrite_wb_0),
	.datad(Mux155),
	.cin(gnd),
	.combout(\reg_file_nxt[31][9]~79_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][9]~79 .lut_mask = 16'hFB00;
defparam \reg_file_nxt[31][9]~79 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N13
dffeas \reg_file[24][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][9] .is_wysiwyg = "true";
defparam \reg_file[24][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N2
cycloneive_lcell_comb \reg_file[16][9]~feeder (
// Equation(s):
// \reg_file[16][9]~feeder_combout  = \reg_file_nxt[31][9]~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][9]~79_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[16][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[16][9]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[16][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N3
dffeas \reg_file[16][9] (
	.clk(!CLK),
	.d(\reg_file[16][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][9] .is_wysiwyg = "true";
defparam \reg_file[16][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N14
cycloneive_lcell_comb \reg_file[20][9]~feeder (
// Equation(s):
// \reg_file[20][9]~feeder_combout  = \reg_file_nxt[31][9]~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][9]~79_combout ),
	.cin(gnd),
	.combout(\reg_file[20][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[20][9]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[20][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N15
dffeas \reg_file[20][9] (
	.clk(!CLK),
	.d(\reg_file[20][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][9] .is_wysiwyg = "true";
defparam \reg_file[20][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N8
cycloneive_lcell_comb \Mux54~4 (
// Equation(s):
// \Mux54~4_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[20][9]~q ))) # (!\prif.imemload_id [18] & (\reg_file[16][9]~q ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[16][9]~q ),
	.datac(\reg_file[20][9]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux54~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~4 .lut_mask = 16'hFA44;
defparam \Mux54~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N3
dffeas \reg_file[28][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][9] .is_wysiwyg = "true";
defparam \reg_file[28][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N10
cycloneive_lcell_comb \Mux54~5 (
// Equation(s):
// \Mux54~5_combout  = (\prif.imemload_id [19] & ((\Mux54~4_combout  & ((\reg_file[28][9]~q ))) # (!\Mux54~4_combout  & (\reg_file[24][9]~q )))) # (!\prif.imemload_id [19] & (((\Mux54~4_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[24][9]~q ),
	.datac(\Mux54~4_combout ),
	.datad(\reg_file[28][9]~q ),
	.cin(gnd),
	.combout(\Mux54~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~5 .lut_mask = 16'hF858;
defparam \Mux54~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N1
dffeas \reg_file[26][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][9] .is_wysiwyg = "true";
defparam \reg_file[26][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N22
cycloneive_lcell_comb \reg_file[30][9]~feeder (
// Equation(s):
// \reg_file[30][9]~feeder_combout  = \reg_file_nxt[31][9]~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][9]~79_combout ),
	.cin(gnd),
	.combout(\reg_file[30][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[30][9]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[30][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N23
dffeas \reg_file[30][9] (
	.clk(!CLK),
	.d(\reg_file[30][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][9] .is_wysiwyg = "true";
defparam \reg_file[30][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N3
dffeas \reg_file[18][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][9] .is_wysiwyg = "true";
defparam \reg_file[18][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N1
dffeas \reg_file[22][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][9] .is_wysiwyg = "true";
defparam \reg_file[22][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N2
cycloneive_lcell_comb \Mux54~2 (
// Equation(s):
// \Mux54~2_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[22][9]~q ))) # (!\prif.imemload_id [18] & (\reg_file[18][9]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][9]~q ),
	.datad(\reg_file[22][9]~q ),
	.cin(gnd),
	.combout(\Mux54~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~2 .lut_mask = 16'hDC98;
defparam \Mux54~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N12
cycloneive_lcell_comb \Mux54~3 (
// Equation(s):
// \Mux54~3_combout  = (\prif.imemload_id [19] & ((\Mux54~2_combout  & ((\reg_file[30][9]~q ))) # (!\Mux54~2_combout  & (\reg_file[26][9]~q )))) # (!\prif.imemload_id [19] & (((\Mux54~2_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[26][9]~q ),
	.datac(\reg_file[30][9]~q ),
	.datad(\Mux54~2_combout ),
	.cin(gnd),
	.combout(\Mux54~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~3 .lut_mask = 16'hF588;
defparam \Mux54~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N12
cycloneive_lcell_comb \Mux54~6 (
// Equation(s):
// \Mux54~6_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\Mux54~3_combout ))) # (!\prif.imemload_id [17] & (\Mux54~5_combout ))))

	.dataa(\Mux54~5_combout ),
	.datab(prifimemload_id_16),
	.datac(prifimemload_id_17),
	.datad(\Mux54~3_combout ),
	.cin(gnd),
	.combout(\Mux54~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~6 .lut_mask = 16'hF2C2;
defparam \Mux54~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N9
dffeas \reg_file[29][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][9] .is_wysiwyg = "true";
defparam \reg_file[29][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y26_N3
dffeas \reg_file[21][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][9] .is_wysiwyg = "true";
defparam \reg_file[21][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y26_N23
dffeas \reg_file[17][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][9] .is_wysiwyg = "true";
defparam \reg_file[17][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y26_N13
dffeas \reg_file[25][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][9] .is_wysiwyg = "true";
defparam \reg_file[25][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N12
cycloneive_lcell_comb \Mux54~0 (
// Equation(s):
// \Mux54~0_combout  = (\prif.imemload_id [19] & (((\reg_file[25][9]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[17][9]~q  & ((!\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[17][9]~q ),
	.datac(\reg_file[25][9]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux54~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~0 .lut_mask = 16'hAAE4;
defparam \Mux54~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N2
cycloneive_lcell_comb \Mux54~1 (
// Equation(s):
// \Mux54~1_combout  = (\prif.imemload_id [18] & ((\Mux54~0_combout  & (\reg_file[29][9]~q )) # (!\Mux54~0_combout  & ((\reg_file[21][9]~q ))))) # (!\prif.imemload_id [18] & (((\Mux54~0_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[29][9]~q ),
	.datac(\reg_file[21][9]~q ),
	.datad(\Mux54~0_combout ),
	.cin(gnd),
	.combout(\Mux54~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~1 .lut_mask = 16'hDDA0;
defparam \Mux54~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N21
dffeas \reg_file[27][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][9] .is_wysiwyg = "true";
defparam \reg_file[27][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N20
cycloneive_lcell_comb \Mux54~7 (
// Equation(s):
// \Mux54~7_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[27][9]~q ))) # (!\prif.imemload_id [19] & (\reg_file[19][9]~q ))))

	.dataa(\reg_file[19][9]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[27][9]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux54~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~7 .lut_mask = 16'hFC22;
defparam \Mux54~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N15
dffeas \reg_file[23][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][9] .is_wysiwyg = "true";
defparam \reg_file[23][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N9
dffeas \reg_file[31][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][9] .is_wysiwyg = "true";
defparam \reg_file[31][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N14
cycloneive_lcell_comb \Mux54~8 (
// Equation(s):
// \Mux54~8_combout  = (\Mux54~7_combout  & (((\reg_file[31][9]~q )) # (!\prif.imemload_id [18]))) # (!\Mux54~7_combout  & (\prif.imemload_id [18] & (\reg_file[23][9]~q )))

	.dataa(\Mux54~7_combout ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[23][9]~q ),
	.datad(\reg_file[31][9]~q ),
	.cin(gnd),
	.combout(\Mux54~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~8 .lut_mask = 16'hEA62;
defparam \Mux54~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N27
dffeas \reg_file[12][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][9] .is_wysiwyg = "true";
defparam \reg_file[12][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N1
dffeas \reg_file[13][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][9] .is_wysiwyg = "true";
defparam \reg_file[13][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N26
cycloneive_lcell_comb \Mux54~17 (
// Equation(s):
// \Mux54~17_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[13][9]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[12][9]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[12][9]~q ),
	.datad(\reg_file[13][9]~q ),
	.cin(gnd),
	.combout(\Mux54~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~17 .lut_mask = 16'hBA98;
defparam \Mux54~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y31_N5
dffeas \reg_file[14][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][9] .is_wysiwyg = "true";
defparam \reg_file[14][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N11
dffeas \reg_file[15][9] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][9]~79_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][9] .is_wysiwyg = "true";
defparam \reg_file[15][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N26
cycloneive_lcell_comb \Mux54~18 (
// Equation(s):
// \Mux54~18_combout  = (\Mux54~17_combout  & (((\reg_file[15][9]~q ) # (!\prif.imemload_id [17])))) # (!\Mux54~17_combout  & (\reg_file[14][9]~q  & (\prif.imemload_id [17])))

	.dataa(\Mux54~17_combout ),
	.datab(\reg_file[14][9]~q ),
	.datac(prifimemload_id_17),
	.datad(\reg_file[15][9]~q ),
	.cin(gnd),
	.combout(\Mux54~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~18 .lut_mask = 16'hEA4A;
defparam \Mux54~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N16
cycloneive_lcell_comb \reg_file[2][9]~feeder (
// Equation(s):
// \reg_file[2][9]~feeder_combout  = \reg_file_nxt[31][9]~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][9]~79_combout ),
	.cin(gnd),
	.combout(\reg_file[2][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][9]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[2][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N17
dffeas \reg_file[2][9] (
	.clk(!CLK),
	.d(\reg_file[2][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][9] .is_wysiwyg = "true";
defparam \reg_file[2][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N15
dffeas \reg_file[1][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][9] .is_wysiwyg = "true";
defparam \reg_file[1][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N25
dffeas \reg_file[3][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][9] .is_wysiwyg = "true";
defparam \reg_file[3][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N24
cycloneive_lcell_comb \Mux54~14 (
// Equation(s):
// \Mux54~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][9]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][9]~q ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[1][9]~q ),
	.datac(\reg_file[3][9]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux54~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~14 .lut_mask = 16'hE400;
defparam \Mux54~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N10
cycloneive_lcell_comb \Mux54~15 (
// Equation(s):
// \Mux54~15_combout  = (\Mux54~14_combout ) # ((!\prif.imemload_id [16] & (\reg_file[2][9]~q  & \prif.imemload_id [17])))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[2][9]~q ),
	.datac(\Mux54~14_combout ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux54~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~15 .lut_mask = 16'hF4F0;
defparam \Mux54~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N4
cycloneive_lcell_comb \reg_file[11][9]~feeder (
// Equation(s):
// \reg_file[11][9]~feeder_combout  = \reg_file_nxt[31][9]~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][9]~79_combout ),
	.cin(gnd),
	.combout(\reg_file[11][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[11][9]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[11][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y31_N5
dffeas \reg_file[11][9] (
	.clk(!CLK),
	.d(\reg_file[11][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][9] .is_wysiwyg = "true";
defparam \reg_file[11][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y31_N9
dffeas \reg_file[9][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][9] .is_wysiwyg = "true";
defparam \reg_file[9][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N26
cycloneive_lcell_comb \Mux54~13 (
// Equation(s):
// \Mux54~13_combout  = (\Mux54~12_combout  & ((\reg_file[11][9]~q ) # ((!\prif.imemload_id [16])))) # (!\Mux54~12_combout  & (((\prif.imemload_id [16] & \reg_file[9][9]~q ))))

	.dataa(\Mux54~12_combout ),
	.datab(\reg_file[11][9]~q ),
	.datac(prifimemload_id_16),
	.datad(\reg_file[9][9]~q ),
	.cin(gnd),
	.combout(\Mux54~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~13 .lut_mask = 16'hDA8A;
defparam \Mux54~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N24
cycloneive_lcell_comb \Mux54~16 (
// Equation(s):
// \Mux54~16_combout  = (\prif.imemload_id [19] & (((\Mux54~13_combout ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\Mux54~15_combout  & ((!\prif.imemload_id [18]))))

	.dataa(\Mux54~15_combout ),
	.datab(prifimemload_id_19),
	.datac(\Mux54~13_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux54~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~16 .lut_mask = 16'hCCE2;
defparam \Mux54~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N30
cycloneive_lcell_comb \reg_file[6][9]~feeder (
// Equation(s):
// \reg_file[6][9]~feeder_combout  = \reg_file_nxt[31][9]~79_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][9]~79_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][9]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][9]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][9]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N31
dffeas \reg_file[6][9] (
	.clk(!CLK),
	.d(\reg_file[6][9]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][9] .is_wysiwyg = "true";
defparam \reg_file[6][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N21
dffeas \reg_file[5][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][9] .is_wysiwyg = "true";
defparam \reg_file[5][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y28_N21
dffeas \reg_file[4][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][9] .is_wysiwyg = "true";
defparam \reg_file[4][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N20
cycloneive_lcell_comb \Mux54~10 (
// Equation(s):
// \Mux54~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][9]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][9]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][9]~q ),
	.datad(\reg_file[4][9]~q ),
	.cin(gnd),
	.combout(\Mux54~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~10 .lut_mask = 16'hB9A8;
defparam \Mux54~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N3
dffeas \reg_file[7][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][9] .is_wysiwyg = "true";
defparam \reg_file[7][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N0
cycloneive_lcell_comb \Mux54~11 (
// Equation(s):
// \Mux54~11_combout  = (\Mux54~10_combout  & (((\reg_file[7][9]~q ) # (!\prif.imemload_id [17])))) # (!\Mux54~10_combout  & (\reg_file[6][9]~q  & ((\prif.imemload_id [17]))))

	.dataa(\reg_file[6][9]~q ),
	.datab(\Mux54~10_combout ),
	.datac(\reg_file[7][9]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux54~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux54~11 .lut_mask = 16'hE2CC;
defparam \Mux54~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N4
cycloneive_lcell_comb \reg_file_nxt[31][6]~80 (
// Equation(s):
// \reg_file_nxt[31][6]~80_combout  = (\Mux158~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Equal8),
	.datac(prifregwrite_wb_0),
	.datad(Mux158),
	.cin(gnd),
	.combout(\reg_file_nxt[31][6]~80_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][6]~80 .lut_mask = 16'hFB00;
defparam \reg_file_nxt[31][6]~80 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N5
dffeas \reg_file[25][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][6] .is_wysiwyg = "true";
defparam \reg_file[25][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N9
dffeas \reg_file[17][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][6] .is_wysiwyg = "true";
defparam \reg_file[17][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N8
cycloneive_lcell_comb \Mux57~0 (
// Equation(s):
// \Mux57~0_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[21][6]~q )) # (!\prif.imemload_id [18] & ((\reg_file[17][6]~q )))))

	.dataa(\reg_file[21][6]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][6]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux57~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~0 .lut_mask = 16'hEE30;
defparam \Mux57~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N0
cycloneive_lcell_comb \reg_file[29][6]~feeder (
// Equation(s):
// \reg_file[29][6]~feeder_combout  = \reg_file_nxt[31][6]~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][6]~80_combout ),
	.cin(gnd),
	.combout(\reg_file[29][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][6]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N1
dffeas \reg_file[29][6] (
	.clk(!CLK),
	.d(\reg_file[29][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][6] .is_wysiwyg = "true";
defparam \reg_file[29][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N8
cycloneive_lcell_comb \Mux57~1 (
// Equation(s):
// \Mux57~1_combout  = (\Mux57~0_combout  & (((\reg_file[29][6]~q ) # (!\prif.imemload_id [19])))) # (!\Mux57~0_combout  & (\reg_file[25][6]~q  & ((\prif.imemload_id [19]))))

	.dataa(\reg_file[25][6]~q ),
	.datab(\Mux57~0_combout ),
	.datac(\reg_file[29][6]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux57~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~1 .lut_mask = 16'hE2CC;
defparam \Mux57~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N9
dffeas \reg_file[23][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][6] .is_wysiwyg = "true";
defparam \reg_file[23][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N25
dffeas \reg_file[19][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][6] .is_wysiwyg = "true";
defparam \reg_file[19][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N8
cycloneive_lcell_comb \Mux57~7 (
// Equation(s):
// \Mux57~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][6]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][6]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][6]~q ),
	.datad(\reg_file[19][6]~q ),
	.cin(gnd),
	.combout(\Mux57~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~7 .lut_mask = 16'hB9A8;
defparam \Mux57~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y27_N3
dffeas \reg_file[31][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][6] .is_wysiwyg = "true";
defparam \reg_file[31][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N8
cycloneive_lcell_comb \reg_file[27][6]~feeder (
// Equation(s):
// \reg_file[27][6]~feeder_combout  = \reg_file_nxt[31][6]~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][6]~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[27][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[27][6]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[27][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N9
dffeas \reg_file[27][6] (
	.clk(!CLK),
	.d(\reg_file[27][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][6] .is_wysiwyg = "true";
defparam \reg_file[27][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N2
cycloneive_lcell_comb \Mux57~8 (
// Equation(s):
// \Mux57~8_combout  = (\prif.imemload_id [19] & ((\Mux57~7_combout  & (\reg_file[31][6]~q )) # (!\Mux57~7_combout  & ((\reg_file[27][6]~q ))))) # (!\prif.imemload_id [19] & (\Mux57~7_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux57~7_combout ),
	.datac(\reg_file[31][6]~q ),
	.datad(\reg_file[27][6]~q ),
	.cin(gnd),
	.combout(\Mux57~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~8 .lut_mask = 16'hE6C4;
defparam \Mux57~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N7
dffeas \reg_file[22][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][6] .is_wysiwyg = "true";
defparam \reg_file[22][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N15
dffeas \reg_file[18][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][6] .is_wysiwyg = "true";
defparam \reg_file[18][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N26
cycloneive_lcell_comb \reg_file[26][6]~feeder (
// Equation(s):
// \reg_file[26][6]~feeder_combout  = \reg_file_nxt[31][6]~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][6]~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[26][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[26][6]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[26][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N27
dffeas \reg_file[26][6] (
	.clk(!CLK),
	.d(\reg_file[26][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][6] .is_wysiwyg = "true";
defparam \reg_file[26][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N14
cycloneive_lcell_comb \Mux57~2 (
// Equation(s):
// \Mux57~2_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[26][6]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & (\reg_file[18][6]~q )))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[18][6]~q ),
	.datad(\reg_file[26][6]~q ),
	.cin(gnd),
	.combout(\Mux57~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~2 .lut_mask = 16'hBA98;
defparam \Mux57~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N14
cycloneive_lcell_comb \Mux57~3 (
// Equation(s):
// \Mux57~3_combout  = (\prif.imemload_id [18] & ((\Mux57~2_combout  & (\reg_file[30][6]~q )) # (!\Mux57~2_combout  & ((\reg_file[22][6]~q ))))) # (!\prif.imemload_id [18] & (((\Mux57~2_combout ))))

	.dataa(\reg_file[30][6]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[22][6]~q ),
	.datad(\Mux57~2_combout ),
	.cin(gnd),
	.combout(\Mux57~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~3 .lut_mask = 16'hBBC0;
defparam \Mux57~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N29
dffeas \reg_file[28][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][6] .is_wysiwyg = "true";
defparam \reg_file[28][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N19
dffeas \reg_file[16][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][6] .is_wysiwyg = "true";
defparam \reg_file[16][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N20
cycloneive_lcell_comb \reg_file[24][6]~feeder (
// Equation(s):
// \reg_file[24][6]~feeder_combout  = \reg_file_nxt[31][6]~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][6]~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[24][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][6]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[24][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N21
dffeas \reg_file[24][6] (
	.clk(!CLK),
	.d(\reg_file[24][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][6] .is_wysiwyg = "true";
defparam \reg_file[24][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N18
cycloneive_lcell_comb \Mux57~4 (
// Equation(s):
// \Mux57~4_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[24][6]~q ))) # (!\prif.imemload_id [19] & (\reg_file[16][6]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[16][6]~q ),
	.datad(\reg_file[24][6]~q ),
	.cin(gnd),
	.combout(\Mux57~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~4 .lut_mask = 16'hDC98;
defparam \Mux57~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N6
cycloneive_lcell_comb \Mux57~5 (
// Equation(s):
// \Mux57~5_combout  = (\Mux57~4_combout  & (((\reg_file[28][6]~q ) # (!\prif.imemload_id [18])))) # (!\Mux57~4_combout  & (\reg_file[20][6]~q  & ((\prif.imemload_id [18]))))

	.dataa(\reg_file[20][6]~q ),
	.datab(\reg_file[28][6]~q ),
	.datac(\Mux57~4_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux57~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~5 .lut_mask = 16'hCAF0;
defparam \Mux57~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N0
cycloneive_lcell_comb \Mux57~6 (
// Equation(s):
// \Mux57~6_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\Mux57~3_combout )) # (!\prif.imemload_id [17] & ((\Mux57~5_combout )))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\Mux57~3_combout ),
	.datad(\Mux57~5_combout ),
	.cin(gnd),
	.combout(\Mux57~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~6 .lut_mask = 16'hD9C8;
defparam \Mux57~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N27
dffeas \reg_file[1][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][6] .is_wysiwyg = "true";
defparam \reg_file[1][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N12
cycloneive_lcell_comb \reg_file[3][6]~feeder (
// Equation(s):
// \reg_file[3][6]~feeder_combout  = \reg_file_nxt[31][6]~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][6]~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[3][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[3][6]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[3][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y28_N13
dffeas \reg_file[3][6] (
	.clk(!CLK),
	.d(\reg_file[3][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][6] .is_wysiwyg = "true";
defparam \reg_file[3][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N26
cycloneive_lcell_comb \Mux57~14 (
// Equation(s):
// \Mux57~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][6]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][6]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[1][6]~q ),
	.datad(\reg_file[3][6]~q ),
	.cin(gnd),
	.combout(\Mux57~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~14 .lut_mask = 16'hA820;
defparam \Mux57~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y28_N21
dffeas \reg_file[2][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][6] .is_wysiwyg = "true";
defparam \reg_file[2][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N20
cycloneive_lcell_comb \Mux57~15 (
// Equation(s):
// \Mux57~15_combout  = (\Mux57~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][6]~q )))

	.dataa(prifimemload_id_16),
	.datab(\Mux57~14_combout ),
	.datac(prifimemload_id_17),
	.datad(\reg_file[2][6]~q ),
	.cin(gnd),
	.combout(\Mux57~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~15 .lut_mask = 16'hDCCC;
defparam \Mux57~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N17
dffeas \reg_file[6][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][6] .is_wysiwyg = "true";
defparam \reg_file[6][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N31
dffeas \reg_file[7][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][6] .is_wysiwyg = "true";
defparam \reg_file[7][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N21
dffeas \reg_file[5][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][6] .is_wysiwyg = "true";
defparam \reg_file[5][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N7
dffeas \reg_file[4][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][6] .is_wysiwyg = "true";
defparam \reg_file[4][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N20
cycloneive_lcell_comb \Mux57~12 (
// Equation(s):
// \Mux57~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][6]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][6]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][6]~q ),
	.datad(\reg_file[4][6]~q ),
	.cin(gnd),
	.combout(\Mux57~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~12 .lut_mask = 16'hB9A8;
defparam \Mux57~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N30
cycloneive_lcell_comb \Mux57~13 (
// Equation(s):
// \Mux57~13_combout  = (\prif.imemload_id [17] & ((\Mux57~12_combout  & ((\reg_file[7][6]~q ))) # (!\Mux57~12_combout  & (\reg_file[6][6]~q )))) # (!\prif.imemload_id [17] & (((\Mux57~12_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][6]~q ),
	.datac(\reg_file[7][6]~q ),
	.datad(\Mux57~12_combout ),
	.cin(gnd),
	.combout(\Mux57~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~13 .lut_mask = 16'hF588;
defparam \Mux57~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N10
cycloneive_lcell_comb \Mux57~16 (
// Equation(s):
// \Mux57~16_combout  = (\prif.imemload_id [18] & (((\Mux57~13_combout ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\Mux57~15_combout  & ((!\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\Mux57~15_combout ),
	.datac(\Mux57~13_combout ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux57~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~16 .lut_mask = 16'hAAE4;
defparam \Mux57~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N9
dffeas \reg_file[9][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][6] .is_wysiwyg = "true";
defparam \reg_file[9][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N3
dffeas \reg_file[11][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][6] .is_wysiwyg = "true";
defparam \reg_file[11][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N9
dffeas \reg_file[10][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][6] .is_wysiwyg = "true";
defparam \reg_file[10][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N11
dffeas \reg_file[8][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][6] .is_wysiwyg = "true";
defparam \reg_file[8][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N10
cycloneive_lcell_comb \Mux57~10 (
// Equation(s):
// \Mux57~10_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[10][6]~q )) # (!\prif.imemload_id [17] & ((\reg_file[8][6]~q )))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[10][6]~q ),
	.datac(\reg_file[8][6]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux57~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~10 .lut_mask = 16'hEE50;
defparam \Mux57~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N2
cycloneive_lcell_comb \Mux57~11 (
// Equation(s):
// \Mux57~11_combout  = (\prif.imemload_id [16] & ((\Mux57~10_combout  & ((\reg_file[11][6]~q ))) # (!\Mux57~10_combout  & (\reg_file[9][6]~q )))) # (!\prif.imemload_id [16] & (((\Mux57~10_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[9][6]~q ),
	.datac(\reg_file[11][6]~q ),
	.datad(\Mux57~10_combout ),
	.cin(gnd),
	.combout(\Mux57~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~11 .lut_mask = 16'hF588;
defparam \Mux57~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N5
dffeas \reg_file[15][6] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][6]~80_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][6] .is_wysiwyg = "true";
defparam \reg_file[15][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N4
cycloneive_lcell_comb \reg_file[14][6]~feeder (
// Equation(s):
// \reg_file[14][6]~feeder_combout  = \reg_file_nxt[31][6]~80_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][6]~80_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[14][6]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][6]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[14][6]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N5
dffeas \reg_file[14][6] (
	.clk(!CLK),
	.d(\reg_file[14][6]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][6] .is_wysiwyg = "true";
defparam \reg_file[14][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N29
dffeas \reg_file[13][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][6] .is_wysiwyg = "true";
defparam \reg_file[13][6] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N3
dffeas \reg_file[12][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][6] .is_wysiwyg = "true";
defparam \reg_file[12][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N28
cycloneive_lcell_comb \Mux57~17 (
// Equation(s):
// \Mux57~17_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[13][6]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[12][6]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[13][6]~q ),
	.datad(\reg_file[12][6]~q ),
	.cin(gnd),
	.combout(\Mux57~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~17 .lut_mask = 16'hB9A8;
defparam \Mux57~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N24
cycloneive_lcell_comb \Mux57~18 (
// Equation(s):
// \Mux57~18_combout  = (\prif.imemload_id [17] & ((\Mux57~17_combout  & (\reg_file[15][6]~q )) # (!\Mux57~17_combout  & ((\reg_file[14][6]~q ))))) # (!\prif.imemload_id [17] & (((\Mux57~17_combout ))))

	.dataa(\reg_file[15][6]~q ),
	.datab(\reg_file[14][6]~q ),
	.datac(prifimemload_id_17),
	.datad(\Mux57~17_combout ),
	.cin(gnd),
	.combout(\Mux57~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux57~18 .lut_mask = 16'hAFC0;
defparam \Mux57~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N30
cycloneive_lcell_comb \reg_file_nxt[31][27]~81 (
// Equation(s):
// \reg_file_nxt[31][27]~81_combout  = (\Mux137~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Mux137),
	.datac(prifregwrite_wb_0),
	.datad(Equal8),
	.cin(gnd),
	.combout(\reg_file_nxt[31][27]~81_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][27]~81 .lut_mask = 16'hC8CC;
defparam \reg_file_nxt[31][27]~81 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N11
dffeas \reg_file[26][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][27] .is_wysiwyg = "true";
defparam \reg_file[26][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N23
dffeas \reg_file[30][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][27] .is_wysiwyg = "true";
defparam \reg_file[30][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N6
cycloneive_lcell_comb \Mux36~3 (
// Equation(s):
// \Mux36~3_combout  = (\Mux36~2_combout  & (((\reg_file[30][27]~q ) # (!\prif.imemload_id [19])))) # (!\Mux36~2_combout  & (\reg_file[26][27]~q  & (\prif.imemload_id [19])))

	.dataa(\Mux36~2_combout ),
	.datab(\reg_file[26][27]~q ),
	.datac(prifimemload_id_19),
	.datad(\reg_file[30][27]~q ),
	.cin(gnd),
	.combout(\Mux36~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~3 .lut_mask = 16'hEA4A;
defparam \Mux36~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N21
dffeas \reg_file[28][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][27] .is_wysiwyg = "true";
defparam \reg_file[28][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N29
dffeas \reg_file[20][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][27] .is_wysiwyg = "true";
defparam \reg_file[20][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N28
cycloneive_lcell_comb \Mux36~4 (
// Equation(s):
// \Mux36~4_combout  = (\prif.imemload_id [18] & (((\reg_file[20][27]~q ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\reg_file[16][27]~q  & ((!\prif.imemload_id [19]))))

	.dataa(\reg_file[16][27]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[20][27]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux36~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~4 .lut_mask = 16'hCCE2;
defparam \Mux36~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N20
cycloneive_lcell_comb \Mux36~5 (
// Equation(s):
// \Mux36~5_combout  = (\prif.imemload_id [19] & ((\Mux36~4_combout  & ((\reg_file[28][27]~q ))) # (!\Mux36~4_combout  & (\reg_file[24][27]~q )))) # (!\prif.imemload_id [19] & (((\Mux36~4_combout ))))

	.dataa(\reg_file[24][27]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[28][27]~q ),
	.datad(\Mux36~4_combout ),
	.cin(gnd),
	.combout(\Mux36~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~5 .lut_mask = 16'hF388;
defparam \Mux36~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N8
cycloneive_lcell_comb \Mux36~6 (
// Equation(s):
// \Mux36~6_combout  = (\prif.imemload_id [17] & ((\Mux36~3_combout ) # ((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (((\Mux36~5_combout  & !\prif.imemload_id [16]))))

	.dataa(prifimemload_id_17),
	.datab(\Mux36~3_combout ),
	.datac(\Mux36~5_combout ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux36~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~6 .lut_mask = 16'hAAD8;
defparam \Mux36~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N6
cycloneive_lcell_comb \reg_file[29][27]~feeder (
// Equation(s):
// \reg_file[29][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][27]~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][27]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N7
dffeas \reg_file[29][27] (
	.clk(!CLK),
	.d(\reg_file[29][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][27] .is_wysiwyg = "true";
defparam \reg_file[29][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y32_N13
dffeas \reg_file[21][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][27] .is_wysiwyg = "true";
defparam \reg_file[21][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N29
dffeas \reg_file[17][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][27] .is_wysiwyg = "true";
defparam \reg_file[17][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N28
cycloneive_lcell_comb \Mux36~0 (
// Equation(s):
// \Mux36~0_combout  = (\prif.imemload_id [19] & ((\reg_file[25][27]~q ) # ((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (((\reg_file[17][27]~q  & !\prif.imemload_id [18]))))

	.dataa(\reg_file[25][27]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][27]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux36~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~0 .lut_mask = 16'hCCB8;
defparam \Mux36~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N12
cycloneive_lcell_comb \Mux36~1 (
// Equation(s):
// \Mux36~1_combout  = (\Mux36~0_combout  & ((\reg_file[29][27]~q ) # ((!\prif.imemload_id [18])))) # (!\Mux36~0_combout  & (((\reg_file[21][27]~q  & \prif.imemload_id [18]))))

	.dataa(\reg_file[29][27]~q ),
	.datab(\reg_file[21][27]~q ),
	.datac(\Mux36~0_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux36~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~1 .lut_mask = 16'hACF0;
defparam \Mux36~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N7
dffeas \reg_file[27][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][27] .is_wysiwyg = "true";
defparam \reg_file[27][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N29
dffeas \reg_file[19][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][27] .is_wysiwyg = "true";
defparam \reg_file[19][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N6
cycloneive_lcell_comb \Mux36~7 (
// Equation(s):
// \Mux36~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][27]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][27]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][27]~q ),
	.datad(\reg_file[19][27]~q ),
	.cin(gnd),
	.combout(\Mux36~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~7 .lut_mask = 16'hD9C8;
defparam \Mux36~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N26
cycloneive_lcell_comb \reg_file[23][27]~feeder (
// Equation(s):
// \reg_file[23][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][27]~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[23][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][27]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[23][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y26_N27
dffeas \reg_file[23][27] (
	.clk(!CLK),
	.d(\reg_file[23][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][27] .is_wysiwyg = "true";
defparam \reg_file[23][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N10
cycloneive_lcell_comb \reg_file[31][27]~feeder (
// Equation(s):
// \reg_file[31][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][27]~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[31][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][27]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[31][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N11
dffeas \reg_file[31][27] (
	.clk(!CLK),
	.d(\reg_file[31][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][27] .is_wysiwyg = "true";
defparam \reg_file[31][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N16
cycloneive_lcell_comb \Mux36~8 (
// Equation(s):
// \Mux36~8_combout  = (\Mux36~7_combout  & (((\reg_file[31][27]~q )) # (!\prif.imemload_id [18]))) # (!\Mux36~7_combout  & (\prif.imemload_id [18] & (\reg_file[23][27]~q )))

	.dataa(\Mux36~7_combout ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[23][27]~q ),
	.datad(\reg_file[31][27]~q ),
	.cin(gnd),
	.combout(\Mux36~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~8 .lut_mask = 16'hEA62;
defparam \Mux36~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N31
dffeas \reg_file[15][27] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][27]~81_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][27] .is_wysiwyg = "true";
defparam \reg_file[15][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N5
dffeas \reg_file[13][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][27] .is_wysiwyg = "true";
defparam \reg_file[13][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N27
dffeas \reg_file[12][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][27] .is_wysiwyg = "true";
defparam \reg_file[12][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N26
cycloneive_lcell_comb \Mux36~17 (
// Equation(s):
// \Mux36~17_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & (\reg_file[13][27]~q )) # (!\prif.imemload_id [16] & ((\reg_file[12][27]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[13][27]~q ),
	.datac(\reg_file[12][27]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux36~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~17 .lut_mask = 16'hEE50;
defparam \Mux36~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N2
cycloneive_lcell_comb \reg_file[14][27]~feeder (
// Equation(s):
// \reg_file[14][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][27]~81_combout ),
	.cin(gnd),
	.combout(\reg_file[14][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][27]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[14][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N3
dffeas \reg_file[14][27] (
	.clk(!CLK),
	.d(\reg_file[14][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][27] .is_wysiwyg = "true";
defparam \reg_file[14][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N12
cycloneive_lcell_comb \Mux36~18 (
// Equation(s):
// \Mux36~18_combout  = (\Mux36~17_combout  & ((\reg_file[15][27]~q ) # ((!\prif.imemload_id [17])))) # (!\Mux36~17_combout  & (((\prif.imemload_id [17] & \reg_file[14][27]~q ))))

	.dataa(\reg_file[15][27]~q ),
	.datab(\Mux36~17_combout ),
	.datac(prifimemload_id_17),
	.datad(\reg_file[14][27]~q ),
	.cin(gnd),
	.combout(\Mux36~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~18 .lut_mask = 16'hBC8C;
defparam \Mux36~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N11
dffeas \reg_file[1][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][27] .is_wysiwyg = "true";
defparam \reg_file[1][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N16
cycloneive_lcell_comb \reg_file[3][27]~feeder (
// Equation(s):
// \reg_file[3][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][27]~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[3][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[3][27]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[3][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N17
dffeas \reg_file[3][27] (
	.clk(!CLK),
	.d(\reg_file[3][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][27] .is_wysiwyg = "true";
defparam \reg_file[3][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N10
cycloneive_lcell_comb \Mux36~14 (
// Equation(s):
// \Mux36~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][27]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][27]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][27]~q ),
	.datad(\reg_file[3][27]~q ),
	.cin(gnd),
	.combout(\Mux36~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~14 .lut_mask = 16'hC840;
defparam \Mux36~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y32_N2
cycloneive_lcell_comb \reg_file[2][27]~feeder (
// Equation(s):
// \reg_file[2][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][27]~81_combout ),
	.cin(gnd),
	.combout(\reg_file[2][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][27]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[2][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y32_N3
dffeas \reg_file[2][27] (
	.clk(!CLK),
	.d(\reg_file[2][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][27] .is_wysiwyg = "true";
defparam \reg_file[2][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N16
cycloneive_lcell_comb \Mux36~15 (
// Equation(s):
// \Mux36~15_combout  = (\Mux36~14_combout ) # ((!\prif.imemload_id [16] & (\reg_file[2][27]~q  & \prif.imemload_id [17])))

	.dataa(prifimemload_id_16),
	.datab(\Mux36~14_combout ),
	.datac(\reg_file[2][27]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux36~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~15 .lut_mask = 16'hDCCC;
defparam \Mux36~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N1
dffeas \reg_file[9][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][27] .is_wysiwyg = "true";
defparam \reg_file[9][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N11
dffeas \reg_file[11][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][27] .is_wysiwyg = "true";
defparam \reg_file[11][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N27
dffeas \reg_file[8][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][27] .is_wysiwyg = "true";
defparam \reg_file[8][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N25
dffeas \reg_file[10][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][27] .is_wysiwyg = "true";
defparam \reg_file[10][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N26
cycloneive_lcell_comb \Mux36~12 (
// Equation(s):
// \Mux36~12_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][27]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][27]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[8][27]~q ),
	.datad(\reg_file[10][27]~q ),
	.cin(gnd),
	.combout(\Mux36~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~12 .lut_mask = 16'hDC98;
defparam \Mux36~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N10
cycloneive_lcell_comb \Mux36~13 (
// Equation(s):
// \Mux36~13_combout  = (\prif.imemload_id [16] & ((\Mux36~12_combout  & ((\reg_file[11][27]~q ))) # (!\Mux36~12_combout  & (\reg_file[9][27]~q )))) # (!\prif.imemload_id [16] & (((\Mux36~12_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[9][27]~q ),
	.datac(\reg_file[11][27]~q ),
	.datad(\Mux36~12_combout ),
	.cin(gnd),
	.combout(\Mux36~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~13 .lut_mask = 16'hF588;
defparam \Mux36~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N30
cycloneive_lcell_comb \Mux36~16 (
// Equation(s):
// \Mux36~16_combout  = (\prif.imemload_id [19] & (((\Mux36~13_combout ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\Mux36~15_combout  & ((!\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\Mux36~15_combout ),
	.datac(\Mux36~13_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux36~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~16 .lut_mask = 16'hAAE4;
defparam \Mux36~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N3
dffeas \reg_file[7][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][27] .is_wysiwyg = "true";
defparam \reg_file[7][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N13
dffeas \reg_file[6][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][27] .is_wysiwyg = "true";
defparam \reg_file[6][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N15
dffeas \reg_file[5][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][27] .is_wysiwyg = "true";
defparam \reg_file[5][27] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N1
dffeas \reg_file[4][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][27] .is_wysiwyg = "true";
defparam \reg_file[4][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N14
cycloneive_lcell_comb \Mux36~10 (
// Equation(s):
// \Mux36~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][27]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][27]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][27]~q ),
	.datad(\reg_file[4][27]~q ),
	.cin(gnd),
	.combout(\Mux36~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~10 .lut_mask = 16'hB9A8;
defparam \Mux36~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N12
cycloneive_lcell_comb \Mux36~11 (
// Equation(s):
// \Mux36~11_combout  = (\prif.imemload_id [17] & ((\Mux36~10_combout  & (\reg_file[7][27]~q )) # (!\Mux36~10_combout  & ((\reg_file[6][27]~q ))))) # (!\prif.imemload_id [17] & (((\Mux36~10_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[7][27]~q ),
	.datac(\reg_file[6][27]~q ),
	.datad(\Mux36~10_combout ),
	.cin(gnd),
	.combout(\Mux36~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux36~11 .lut_mask = 16'hDDA0;
defparam \Mux36~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N20
cycloneive_lcell_comb \reg_file_nxt[31][23]~82 (
// Equation(s):
// \reg_file_nxt[31][23]~82_combout  = (\Mux141~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Equal8),
	.datac(prifregwrite_wb_0),
	.datad(Mux141),
	.cin(gnd),
	.combout(\reg_file_nxt[31][23]~82_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][23]~82 .lut_mask = 16'hFB00;
defparam \reg_file_nxt[31][23]~82 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N20
cycloneive_lcell_comb \reg_file[21][23]~feeder (
// Equation(s):
// \reg_file[21][23]~feeder_combout  = \reg_file_nxt[31][23]~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][23]~82_combout ),
	.cin(gnd),
	.combout(\reg_file[21][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][23]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[21][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y32_N21
dffeas \reg_file[21][23] (
	.clk(!CLK),
	.d(\reg_file[21][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][23] .is_wysiwyg = "true";
defparam \reg_file[21][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N15
dffeas \reg_file[25][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][23] .is_wysiwyg = "true";
defparam \reg_file[25][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N14
cycloneive_lcell_comb \Mux40~0 (
// Equation(s):
// \Mux40~0_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[25][23]~q ))) # (!\prif.imemload_id [19] & (\reg_file[17][23]~q ))))

	.dataa(\reg_file[17][23]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[25][23]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux40~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~0 .lut_mask = 16'hFC22;
defparam \Mux40~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N10
cycloneive_lcell_comb \reg_file[29][23]~feeder (
// Equation(s):
// \reg_file[29][23]~feeder_combout  = \reg_file_nxt[31][23]~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][23]~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][23]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N11
dffeas \reg_file[29][23] (
	.clk(!CLK),
	.d(\reg_file[29][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][23] .is_wysiwyg = "true";
defparam \reg_file[29][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N22
cycloneive_lcell_comb \Mux40~1 (
// Equation(s):
// \Mux40~1_combout  = (\prif.imemload_id [18] & ((\Mux40~0_combout  & ((\reg_file[29][23]~q ))) # (!\Mux40~0_combout  & (\reg_file[21][23]~q )))) # (!\prif.imemload_id [18] & (((\Mux40~0_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[21][23]~q ),
	.datac(\Mux40~0_combout ),
	.datad(\reg_file[29][23]~q ),
	.cin(gnd),
	.combout(\Mux40~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~1 .lut_mask = 16'hF858;
defparam \Mux40~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N31
dffeas \reg_file[18][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][23] .is_wysiwyg = "true";
defparam \reg_file[18][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y30_N9
dffeas \reg_file[22][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][23] .is_wysiwyg = "true";
defparam \reg_file[22][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N8
cycloneive_lcell_comb \Mux40~2 (
// Equation(s):
// \Mux40~2_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[22][23]~q ))) # (!\prif.imemload_id [18] & (\reg_file[18][23]~q ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[18][23]~q ),
	.datac(\reg_file[22][23]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux40~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~2 .lut_mask = 16'hFA44;
defparam \Mux40~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N11
dffeas \reg_file[30][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][23] .is_wysiwyg = "true";
defparam \reg_file[30][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N28
cycloneive_lcell_comb \reg_file[26][23]~feeder (
// Equation(s):
// \reg_file[26][23]~feeder_combout  = \reg_file_nxt[31][23]~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][23]~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[26][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[26][23]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[26][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N29
dffeas \reg_file[26][23] (
	.clk(!CLK),
	.d(\reg_file[26][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][23] .is_wysiwyg = "true";
defparam \reg_file[26][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N10
cycloneive_lcell_comb \Mux40~3 (
// Equation(s):
// \Mux40~3_combout  = (\prif.imemload_id [19] & ((\Mux40~2_combout  & (\reg_file[30][23]~q )) # (!\Mux40~2_combout  & ((\reg_file[26][23]~q ))))) # (!\prif.imemload_id [19] & (\Mux40~2_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux40~2_combout ),
	.datac(\reg_file[30][23]~q ),
	.datad(\reg_file[26][23]~q ),
	.cin(gnd),
	.combout(\Mux40~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~3 .lut_mask = 16'hE6C4;
defparam \Mux40~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N17
dffeas \reg_file[28][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][23] .is_wysiwyg = "true";
defparam \reg_file[28][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y34_N19
dffeas \reg_file[24][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][23] .is_wysiwyg = "true";
defparam \reg_file[24][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N18
cycloneive_lcell_comb \Mux40~5 (
// Equation(s):
// \Mux40~5_combout  = (\Mux40~4_combout  & ((\reg_file[28][23]~q ) # ((!\prif.imemload_id [19])))) # (!\Mux40~4_combout  & (((\reg_file[24][23]~q  & \prif.imemload_id [19]))))

	.dataa(\Mux40~4_combout ),
	.datab(\reg_file[28][23]~q ),
	.datac(\reg_file[24][23]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux40~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~5 .lut_mask = 16'hD8AA;
defparam \Mux40~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N4
cycloneive_lcell_comb \Mux40~6 (
// Equation(s):
// \Mux40~6_combout  = (\prif.imemload_id [17] & ((\Mux40~3_combout ) # ((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (((!\prif.imemload_id [16] & \Mux40~5_combout ))))

	.dataa(\Mux40~3_combout ),
	.datab(prifimemload_id_17),
	.datac(prifimemload_id_16),
	.datad(\Mux40~5_combout ),
	.cin(gnd),
	.combout(\Mux40~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~6 .lut_mask = 16'hCBC8;
defparam \Mux40~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N27
dffeas \reg_file[27][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][23] .is_wysiwyg = "true";
defparam \reg_file[27][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N7
dffeas \reg_file[19][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][23] .is_wysiwyg = "true";
defparam \reg_file[19][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N26
cycloneive_lcell_comb \Mux40~7 (
// Equation(s):
// \Mux40~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][23]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][23]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][23]~q ),
	.datad(\reg_file[19][23]~q ),
	.cin(gnd),
	.combout(\Mux40~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~7 .lut_mask = 16'hD9C8;
defparam \Mux40~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N1
dffeas \reg_file[23][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][23] .is_wysiwyg = "true";
defparam \reg_file[23][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N16
cycloneive_lcell_comb \reg_file[31][23]~feeder (
// Equation(s):
// \reg_file[31][23]~feeder_combout  = \reg_file_nxt[31][23]~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][23]~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[31][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][23]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[31][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N17
dffeas \reg_file[31][23] (
	.clk(!CLK),
	.d(\reg_file[31][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][23] .is_wysiwyg = "true";
defparam \reg_file[31][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N0
cycloneive_lcell_comb \Mux40~8 (
// Equation(s):
// \Mux40~8_combout  = (\Mux40~7_combout  & (((\reg_file[31][23]~q )) # (!\prif.imemload_id [18]))) # (!\Mux40~7_combout  & (\prif.imemload_id [18] & (\reg_file[23][23]~q )))

	.dataa(\Mux40~7_combout ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[23][23]~q ),
	.datad(\reg_file[31][23]~q ),
	.cin(gnd),
	.combout(\Mux40~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~8 .lut_mask = 16'hEA62;
defparam \Mux40~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N27
dffeas \reg_file[14][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][23] .is_wysiwyg = "true";
defparam \reg_file[14][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N21
dffeas \reg_file[15][23] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][23]~82_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][23] .is_wysiwyg = "true";
defparam \reg_file[15][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N19
dffeas \reg_file[12][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][23] .is_wysiwyg = "true";
defparam \reg_file[12][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N1
dffeas \reg_file[13][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][23] .is_wysiwyg = "true";
defparam \reg_file[13][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N18
cycloneive_lcell_comb \Mux40~17 (
// Equation(s):
// \Mux40~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][23]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][23]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][23]~q ),
	.datad(\reg_file[13][23]~q ),
	.cin(gnd),
	.combout(\Mux40~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~17 .lut_mask = 16'hDC98;
defparam \Mux40~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N16
cycloneive_lcell_comb \Mux40~18 (
// Equation(s):
// \Mux40~18_combout  = (\prif.imemload_id [17] & ((\Mux40~17_combout  & ((\reg_file[15][23]~q ))) # (!\Mux40~17_combout  & (\reg_file[14][23]~q )))) # (!\prif.imemload_id [17] & (((\Mux40~17_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[14][23]~q ),
	.datac(\reg_file[15][23]~q ),
	.datad(\Mux40~17_combout ),
	.cin(gnd),
	.combout(\Mux40~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~18 .lut_mask = 16'hF588;
defparam \Mux40~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N8
cycloneive_lcell_comb \reg_file[6][23]~feeder (
// Equation(s):
// \reg_file[6][23]~feeder_combout  = \reg_file_nxt[31][23]~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][23]~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][23]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N9
dffeas \reg_file[6][23] (
	.clk(!CLK),
	.d(\reg_file[6][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][23] .is_wysiwyg = "true";
defparam \reg_file[6][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N4
cycloneive_lcell_comb \reg_file[7][23]~feeder (
// Equation(s):
// \reg_file[7][23]~feeder_combout  = \reg_file_nxt[31][23]~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][23]~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[7][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[7][23]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[7][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N5
dffeas \reg_file[7][23] (
	.clk(!CLK),
	.d(\reg_file[7][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][23] .is_wysiwyg = "true";
defparam \reg_file[7][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N23
dffeas \reg_file[5][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][23] .is_wysiwyg = "true";
defparam \reg_file[5][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N17
dffeas \reg_file[4][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][23] .is_wysiwyg = "true";
defparam \reg_file[4][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N22
cycloneive_lcell_comb \Mux40~10 (
// Equation(s):
// \Mux40~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][23]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][23]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][23]~q ),
	.datad(\reg_file[4][23]~q ),
	.cin(gnd),
	.combout(\Mux40~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~10 .lut_mask = 16'hB9A8;
defparam \Mux40~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N26
cycloneive_lcell_comb \Mux40~11 (
// Equation(s):
// \Mux40~11_combout  = (\prif.imemload_id [17] & ((\Mux40~10_combout  & ((\reg_file[7][23]~q ))) # (!\Mux40~10_combout  & (\reg_file[6][23]~q )))) # (!\prif.imemload_id [17] & (((\Mux40~10_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][23]~q ),
	.datac(\reg_file[7][23]~q ),
	.datad(\Mux40~10_combout ),
	.cin(gnd),
	.combout(\Mux40~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~11 .lut_mask = 16'hF588;
defparam \Mux40~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N15
dffeas \reg_file[8][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][23] .is_wysiwyg = "true";
defparam \reg_file[8][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N21
dffeas \reg_file[10][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][23] .is_wysiwyg = "true";
defparam \reg_file[10][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N14
cycloneive_lcell_comb \Mux40~12 (
// Equation(s):
// \Mux40~12_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][23]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][23]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[8][23]~q ),
	.datad(\reg_file[10][23]~q ),
	.cin(gnd),
	.combout(\Mux40~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~12 .lut_mask = 16'hDC98;
defparam \Mux40~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N31
dffeas \reg_file[11][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][23] .is_wysiwyg = "true";
defparam \reg_file[11][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N30
cycloneive_lcell_comb \Mux40~13 (
// Equation(s):
// \Mux40~13_combout  = (\Mux40~12_combout  & (((\reg_file[11][23]~q ) # (!\prif.imemload_id [16])))) # (!\Mux40~12_combout  & (\reg_file[9][23]~q  & ((\prif.imemload_id [16]))))

	.dataa(\reg_file[9][23]~q ),
	.datab(\Mux40~12_combout ),
	.datac(\reg_file[11][23]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux40~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~13 .lut_mask = 16'hE2CC;
defparam \Mux40~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N6
cycloneive_lcell_comb \reg_file[2][23]~feeder (
// Equation(s):
// \reg_file[2][23]~feeder_combout  = \reg_file_nxt[31][23]~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][23]~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[2][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][23]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[2][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N7
dffeas \reg_file[2][23] (
	.clk(!CLK),
	.d(\reg_file[2][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][23] .is_wysiwyg = "true";
defparam \reg_file[2][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N25
dffeas \reg_file[3][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][23] .is_wysiwyg = "true";
defparam \reg_file[3][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N27
dffeas \reg_file[1][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][23] .is_wysiwyg = "true";
defparam \reg_file[1][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N26
cycloneive_lcell_comb \Mux40~14 (
// Equation(s):
// \Mux40~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][23]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][23]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[3][23]~q ),
	.datac(\reg_file[1][23]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux40~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~14 .lut_mask = 16'hD800;
defparam \Mux40~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N24
cycloneive_lcell_comb \Mux40~15 (
// Equation(s):
// \Mux40~15_combout  = (\Mux40~14_combout ) # ((\prif.imemload_id [17] & (\reg_file[2][23]~q  & !\prif.imemload_id [16])))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[2][23]~q ),
	.datac(prifimemload_id_16),
	.datad(\Mux40~14_combout ),
	.cin(gnd),
	.combout(\Mux40~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~15 .lut_mask = 16'hFF08;
defparam \Mux40~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N10
cycloneive_lcell_comb \Mux40~16 (
// Equation(s):
// \Mux40~16_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\Mux40~13_combout )) # (!\prif.imemload_id [19] & ((\Mux40~15_combout )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux40~13_combout ),
	.datad(\Mux40~15_combout ),
	.cin(gnd),
	.combout(\Mux40~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux40~16 .lut_mask = 16'hD9C8;
defparam \Mux40~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N6
cycloneive_lcell_comb \reg_file_nxt[31][18]~83 (
// Equation(s):
// \reg_file_nxt[31][18]~83_combout  = (\Mux146~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Equal8),
	.datac(prifregwrite_wb_0),
	.datad(Mux146),
	.cin(gnd),
	.combout(\reg_file_nxt[31][18]~83_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][18]~83 .lut_mask = 16'hFB00;
defparam \reg_file_nxt[31][18]~83 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N26
cycloneive_lcell_comb \reg_file[30][18]~feeder (
// Equation(s):
// \reg_file[30][18]~feeder_combout  = \reg_file_nxt[31][18]~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][18]~83_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[30][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[30][18]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[30][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N27
dffeas \reg_file[30][18] (
	.clk(!CLK),
	.d(\reg_file[30][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][18] .is_wysiwyg = "true";
defparam \reg_file[30][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N12
cycloneive_lcell_comb \reg_file[22][18]~feeder (
// Equation(s):
// \reg_file[22][18]~feeder_combout  = \reg_file_nxt[31][18]~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][18]~83_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[22][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][18]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[22][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N13
dffeas \reg_file[22][18] (
	.clk(!CLK),
	.d(\reg_file[22][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][18] .is_wysiwyg = "true";
defparam \reg_file[22][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N15
dffeas \reg_file[18][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][18] .is_wysiwyg = "true";
defparam \reg_file[18][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N19
dffeas \reg_file[26][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][18] .is_wysiwyg = "true";
defparam \reg_file[26][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N18
cycloneive_lcell_comb \Mux45~2 (
// Equation(s):
// \Mux45~2_combout  = (\prif.imemload_id [19] & (((\reg_file[26][18]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[18][18]~q  & ((!\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[18][18]~q ),
	.datac(\reg_file[26][18]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux45~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~2 .lut_mask = 16'hAAE4;
defparam \Mux45~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N8
cycloneive_lcell_comb \Mux45~3 (
// Equation(s):
// \Mux45~3_combout  = (\prif.imemload_id [18] & ((\Mux45~2_combout  & (\reg_file[30][18]~q )) # (!\Mux45~2_combout  & ((\reg_file[22][18]~q ))))) # (!\prif.imemload_id [18] & (((\Mux45~2_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[30][18]~q ),
	.datac(\reg_file[22][18]~q ),
	.datad(\Mux45~2_combout ),
	.cin(gnd),
	.combout(\Mux45~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~3 .lut_mask = 16'hDDA0;
defparam \Mux45~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N9
dffeas \reg_file[20][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][18] .is_wysiwyg = "true";
defparam \reg_file[20][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N3
dffeas \reg_file[28][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][18] .is_wysiwyg = "true";
defparam \reg_file[28][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N8
cycloneive_lcell_comb \Mux45~5 (
// Equation(s):
// \Mux45~5_combout  = (\Mux45~4_combout  & (((\reg_file[28][18]~q )) # (!\prif.imemload_id [18]))) # (!\Mux45~4_combout  & (\prif.imemload_id [18] & (\reg_file[20][18]~q )))

	.dataa(\Mux45~4_combout ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[20][18]~q ),
	.datad(\reg_file[28][18]~q ),
	.cin(gnd),
	.combout(\Mux45~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~5 .lut_mask = 16'hEA62;
defparam \Mux45~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N26
cycloneive_lcell_comb \Mux45~6 (
// Equation(s):
// \Mux45~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux45~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & ((\Mux45~5_combout ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux45~3_combout ),
	.datad(\Mux45~5_combout ),
	.cin(gnd),
	.combout(\Mux45~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~6 .lut_mask = 16'hB9A8;
defparam \Mux45~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N15
dffeas \reg_file[23][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][18] .is_wysiwyg = "true";
defparam \reg_file[23][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N9
dffeas \reg_file[19][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][18] .is_wysiwyg = "true";
defparam \reg_file[19][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N14
cycloneive_lcell_comb \Mux45~7 (
// Equation(s):
// \Mux45~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][18]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][18]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][18]~q ),
	.datad(\reg_file[19][18]~q ),
	.cin(gnd),
	.combout(\Mux45~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~7 .lut_mask = 16'hB9A8;
defparam \Mux45~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N17
dffeas \reg_file[27][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][18] .is_wysiwyg = "true";
defparam \reg_file[27][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N15
dffeas \reg_file[31][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][18] .is_wysiwyg = "true";
defparam \reg_file[31][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N16
cycloneive_lcell_comb \Mux45~8 (
// Equation(s):
// \Mux45~8_combout  = (\prif.imemload_id [19] & ((\Mux45~7_combout  & ((\reg_file[31][18]~q ))) # (!\Mux45~7_combout  & (\reg_file[27][18]~q )))) # (!\prif.imemload_id [19] & (\Mux45~7_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux45~7_combout ),
	.datac(\reg_file[27][18]~q ),
	.datad(\reg_file[31][18]~q ),
	.cin(gnd),
	.combout(\Mux45~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~8 .lut_mask = 16'hEC64;
defparam \Mux45~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N29
dffeas \reg_file[25][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][18] .is_wysiwyg = "true";
defparam \reg_file[25][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N18
cycloneive_lcell_comb \reg_file[29][18]~feeder (
// Equation(s):
// \reg_file[29][18]~feeder_combout  = \reg_file_nxt[31][18]~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][18]~83_combout ),
	.cin(gnd),
	.combout(\reg_file[29][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][18]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N19
dffeas \reg_file[29][18] (
	.clk(!CLK),
	.d(\reg_file[29][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][18] .is_wysiwyg = "true";
defparam \reg_file[29][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N31
dffeas \reg_file[17][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][18] .is_wysiwyg = "true";
defparam \reg_file[17][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N2
cycloneive_lcell_comb \reg_file[21][18]~feeder (
// Equation(s):
// \reg_file[21][18]~feeder_combout  = \reg_file_nxt[31][18]~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][18]~83_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[21][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][18]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[21][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N3
dffeas \reg_file[21][18] (
	.clk(!CLK),
	.d(\reg_file[21][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][18] .is_wysiwyg = "true";
defparam \reg_file[21][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N30
cycloneive_lcell_comb \Mux45~0 (
// Equation(s):
// \Mux45~0_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[21][18]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & (\reg_file[17][18]~q )))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][18]~q ),
	.datad(\reg_file[21][18]~q ),
	.cin(gnd),
	.combout(\Mux45~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~0 .lut_mask = 16'hBA98;
defparam \Mux45~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N16
cycloneive_lcell_comb \Mux45~1 (
// Equation(s):
// \Mux45~1_combout  = (\Mux45~0_combout  & (((\reg_file[29][18]~q ) # (!\prif.imemload_id [19])))) # (!\Mux45~0_combout  & (\reg_file[25][18]~q  & ((\prif.imemload_id [19]))))

	.dataa(\reg_file[25][18]~q ),
	.datab(\reg_file[29][18]~q ),
	.datac(\Mux45~0_combout ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux45~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~1 .lut_mask = 16'hCAF0;
defparam \Mux45~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N27
dffeas \reg_file[7][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][18] .is_wysiwyg = "true";
defparam \reg_file[7][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N21
dffeas \reg_file[6][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][18] .is_wysiwyg = "true";
defparam \reg_file[6][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N26
cycloneive_lcell_comb \Mux45~13 (
// Equation(s):
// \Mux45~13_combout  = (\Mux45~12_combout  & (((\reg_file[7][18]~q )) # (!\prif.imemload_id [17]))) # (!\Mux45~12_combout  & (\prif.imemload_id [17] & ((\reg_file[6][18]~q ))))

	.dataa(\Mux45~12_combout ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[7][18]~q ),
	.datad(\reg_file[6][18]~q ),
	.cin(gnd),
	.combout(\Mux45~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~13 .lut_mask = 16'hE6A2;
defparam \Mux45~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N21
dffeas \reg_file[1][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][18] .is_wysiwyg = "true";
defparam \reg_file[1][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N20
cycloneive_lcell_comb \Mux45~14 (
// Equation(s):
// \Mux45~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][18]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][18]~q )))))

	.dataa(\reg_file[3][18]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][18]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux45~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~14 .lut_mask = 16'h88C0;
defparam \Mux45~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N6
cycloneive_lcell_comb \Mux45~15 (
// Equation(s):
// \Mux45~15_combout  = (\Mux45~14_combout ) # ((\reg_file[2][18]~q  & (!\prif.imemload_id [16] & \prif.imemload_id [17])))

	.dataa(\reg_file[2][18]~q ),
	.datab(prifimemload_id_16),
	.datac(\Mux45~14_combout ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux45~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~15 .lut_mask = 16'hF2F0;
defparam \Mux45~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N12
cycloneive_lcell_comb \Mux45~16 (
// Equation(s):
// \Mux45~16_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\Mux45~13_combout )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\Mux45~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux45~13_combout ),
	.datad(\Mux45~15_combout ),
	.cin(gnd),
	.combout(\Mux45~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~16 .lut_mask = 16'hB9A8;
defparam \Mux45~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N8
cycloneive_lcell_comb \reg_file[14][18]~feeder (
// Equation(s):
// \reg_file[14][18]~feeder_combout  = \reg_file_nxt[31][18]~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][18]~83_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[14][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][18]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[14][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N9
dffeas \reg_file[14][18] (
	.clk(!CLK),
	.d(\reg_file[14][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][18] .is_wysiwyg = "true";
defparam \reg_file[14][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y29_N7
dffeas \reg_file[15][18] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][18]~83_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][18] .is_wysiwyg = "true";
defparam \reg_file[15][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N13
dffeas \reg_file[13][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][18] .is_wysiwyg = "true";
defparam \reg_file[13][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N12
cycloneive_lcell_comb \Mux45~17 (
// Equation(s):
// \Mux45~17_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][18]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][18]~q ))))

	.dataa(\reg_file[12][18]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[13][18]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux45~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~17 .lut_mask = 16'hFC22;
defparam \Mux45~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N22
cycloneive_lcell_comb \Mux45~18 (
// Equation(s):
// \Mux45~18_combout  = (\prif.imemload_id [17] & ((\Mux45~17_combout  & ((\reg_file[15][18]~q ))) # (!\Mux45~17_combout  & (\reg_file[14][18]~q )))) # (!\prif.imemload_id [17] & (((\Mux45~17_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[14][18]~q ),
	.datac(\reg_file[15][18]~q ),
	.datad(\Mux45~17_combout ),
	.cin(gnd),
	.combout(\Mux45~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~18 .lut_mask = 16'hF588;
defparam \Mux45~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N28
cycloneive_lcell_comb \reg_file[11][18]~feeder (
// Equation(s):
// \reg_file[11][18]~feeder_combout  = \reg_file_nxt[31][18]~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][18]~83_combout ),
	.cin(gnd),
	.combout(\reg_file[11][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[11][18]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[11][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N29
dffeas \reg_file[11][18] (
	.clk(!CLK),
	.d(\reg_file[11][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][18] .is_wysiwyg = "true";
defparam \reg_file[11][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N17
dffeas \reg_file[9][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][18] .is_wysiwyg = "true";
defparam \reg_file[9][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N19
dffeas \reg_file[8][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][18] .is_wysiwyg = "true";
defparam \reg_file[8][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N1
dffeas \reg_file[10][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][18] .is_wysiwyg = "true";
defparam \reg_file[10][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N0
cycloneive_lcell_comb \Mux45~10 (
// Equation(s):
// \Mux45~10_combout  = (\prif.imemload_id [17] & (((\reg_file[10][18]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][18]~q  & ((!\prif.imemload_id [16]))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[8][18]~q ),
	.datac(\reg_file[10][18]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux45~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~10 .lut_mask = 16'hAAE4;
defparam \Mux45~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N16
cycloneive_lcell_comb \Mux45~11 (
// Equation(s):
// \Mux45~11_combout  = (\prif.imemload_id [16] & ((\Mux45~10_combout  & (\reg_file[11][18]~q )) # (!\Mux45~10_combout  & ((\reg_file[9][18]~q ))))) # (!\prif.imemload_id [16] & (((\Mux45~10_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[11][18]~q ),
	.datac(\reg_file[9][18]~q ),
	.datad(\Mux45~10_combout ),
	.cin(gnd),
	.combout(\Mux45~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux45~11 .lut_mask = 16'hDDA0;
defparam \Mux45~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N8
cycloneive_lcell_comb \reg_file_nxt[31][24]~84 (
// Equation(s):
// \reg_file_nxt[31][24]~84_combout  = (\Mux140~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(Equal8),
	.datac(prifregwrite_wb_0),
	.datad(Mux140),
	.cin(gnd),
	.combout(\reg_file_nxt[31][24]~84_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][24]~84 .lut_mask = 16'hFB00;
defparam \reg_file_nxt[31][24]~84 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N22
cycloneive_lcell_comb \reg_file[29][24]~feeder (
// Equation(s):
// \reg_file[29][24]~feeder_combout  = \reg_file_nxt[31][24]~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][24]~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][24]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N23
dffeas \reg_file[29][24] (
	.clk(!CLK),
	.d(\reg_file[29][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][24] .is_wysiwyg = "true";
defparam \reg_file[29][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N9
dffeas \reg_file[25][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][24] .is_wysiwyg = "true";
defparam \reg_file[25][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N1
dffeas \reg_file[17][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][24] .is_wysiwyg = "true";
defparam \reg_file[17][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N28
cycloneive_lcell_comb \reg_file[21][24]~feeder (
// Equation(s):
// \reg_file[21][24]~feeder_combout  = \reg_file_nxt[31][24]~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][24]~84_combout ),
	.cin(gnd),
	.combout(\reg_file[21][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][24]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[21][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N29
dffeas \reg_file[21][24] (
	.clk(!CLK),
	.d(\reg_file[21][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][24] .is_wysiwyg = "true";
defparam \reg_file[21][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N0
cycloneive_lcell_comb \Mux39~0 (
// Equation(s):
// \Mux39~0_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[21][24]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & (\reg_file[17][24]~q )))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][24]~q ),
	.datad(\reg_file[21][24]~q ),
	.cin(gnd),
	.combout(\Mux39~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~0 .lut_mask = 16'hBA98;
defparam \Mux39~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N10
cycloneive_lcell_comb \Mux39~1 (
// Equation(s):
// \Mux39~1_combout  = (\prif.imemload_id [19] & ((\Mux39~0_combout  & (\reg_file[29][24]~q )) # (!\Mux39~0_combout  & ((\reg_file[25][24]~q ))))) # (!\prif.imemload_id [19] & (((\Mux39~0_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[29][24]~q ),
	.datac(\reg_file[25][24]~q ),
	.datad(\Mux39~0_combout ),
	.cin(gnd),
	.combout(\Mux39~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~1 .lut_mask = 16'hDDA0;
defparam \Mux39~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N7
dffeas \reg_file[28][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][24] .is_wysiwyg = "true";
defparam \reg_file[28][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N25
dffeas \reg_file[16][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][24] .is_wysiwyg = "true";
defparam \reg_file[16][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N24
cycloneive_lcell_comb \Mux39~4 (
// Equation(s):
// \Mux39~4_combout  = (\prif.imemload_id [19] & ((\reg_file[24][24]~q ) # ((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (((\reg_file[16][24]~q  & !\prif.imemload_id [18]))))

	.dataa(\reg_file[24][24]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[16][24]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux39~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~4 .lut_mask = 16'hCCB8;
defparam \Mux39~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N26
cycloneive_lcell_comb \Mux39~5 (
// Equation(s):
// \Mux39~5_combout  = (\prif.imemload_id [18] & ((\Mux39~4_combout  & ((\reg_file[28][24]~q ))) # (!\Mux39~4_combout  & (\reg_file[20][24]~q )))) # (!\prif.imemload_id [18] & (((\Mux39~4_combout ))))

	.dataa(\reg_file[20][24]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[28][24]~q ),
	.datad(\Mux39~4_combout ),
	.cin(gnd),
	.combout(\Mux39~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~5 .lut_mask = 16'hF388;
defparam \Mux39~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N25
dffeas \reg_file[26][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][24] .is_wysiwyg = "true";
defparam \reg_file[26][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N24
cycloneive_lcell_comb \Mux39~2 (
// Equation(s):
// \Mux39~2_combout  = (\prif.imemload_id [19] & (((\reg_file[26][24]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[18][24]~q  & ((!\prif.imemload_id [18]))))

	.dataa(\reg_file[18][24]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[26][24]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux39~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~2 .lut_mask = 16'hCCE2;
defparam \Mux39~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N25
dffeas \reg_file[22][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][24] .is_wysiwyg = "true";
defparam \reg_file[22][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N24
cycloneive_lcell_comb \Mux39~3 (
// Equation(s):
// \Mux39~3_combout  = (\Mux39~2_combout  & ((\reg_file[30][24]~q ) # ((!\prif.imemload_id [18])))) # (!\Mux39~2_combout  & (((\reg_file[22][24]~q  & \prif.imemload_id [18]))))

	.dataa(\reg_file[30][24]~q ),
	.datab(\Mux39~2_combout ),
	.datac(\reg_file[22][24]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux39~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~3 .lut_mask = 16'hB8CC;
defparam \Mux39~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N12
cycloneive_lcell_comb \Mux39~6 (
// Equation(s):
// \Mux39~6_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16]) # (\Mux39~3_combout )))) # (!\prif.imemload_id [17] & (\Mux39~5_combout  & (!\prif.imemload_id [16])))

	.dataa(prifimemload_id_17),
	.datab(\Mux39~5_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux39~3_combout ),
	.cin(gnd),
	.combout(\Mux39~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~6 .lut_mask = 16'hAEA4;
defparam \Mux39~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N14
cycloneive_lcell_comb \reg_file[31][24]~feeder (
// Equation(s):
// \reg_file[31][24]~feeder_combout  = \reg_file_nxt[31][24]~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][24]~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[31][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][24]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[31][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N15
dffeas \reg_file[31][24] (
	.clk(!CLK),
	.d(\reg_file[31][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][24] .is_wysiwyg = "true";
defparam \reg_file[31][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N17
dffeas \reg_file[27][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][24] .is_wysiwyg = "true";
defparam \reg_file[27][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N29
dffeas \reg_file[23][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][24] .is_wysiwyg = "true";
defparam \reg_file[23][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N19
dffeas \reg_file[19][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][24] .is_wysiwyg = "true";
defparam \reg_file[19][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N28
cycloneive_lcell_comb \Mux39~7 (
// Equation(s):
// \Mux39~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][24]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][24]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][24]~q ),
	.datad(\reg_file[19][24]~q ),
	.cin(gnd),
	.combout(\Mux39~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~7 .lut_mask = 16'hB9A8;
defparam \Mux39~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N16
cycloneive_lcell_comb \Mux39~8 (
// Equation(s):
// \Mux39~8_combout  = (\prif.imemload_id [19] & ((\Mux39~7_combout  & (\reg_file[31][24]~q )) # (!\Mux39~7_combout  & ((\reg_file[27][24]~q ))))) # (!\prif.imemload_id [19] & (((\Mux39~7_combout ))))

	.dataa(\reg_file[31][24]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][24]~q ),
	.datad(\Mux39~7_combout ),
	.cin(gnd),
	.combout(\Mux39~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~8 .lut_mask = 16'hBBC0;
defparam \Mux39~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N5
dffeas \reg_file[6][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][24] .is_wysiwyg = "true";
defparam \reg_file[6][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N11
dffeas \reg_file[7][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][24] .is_wysiwyg = "true";
defparam \reg_file[7][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N27
dffeas \reg_file[4][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][24] .is_wysiwyg = "true";
defparam \reg_file[4][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N17
dffeas \reg_file[5][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][24] .is_wysiwyg = "true";
defparam \reg_file[5][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N26
cycloneive_lcell_comb \Mux39~12 (
// Equation(s):
// \Mux39~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][24]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][24]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][24]~q ),
	.datad(\reg_file[5][24]~q ),
	.cin(gnd),
	.combout(\Mux39~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~12 .lut_mask = 16'hBA98;
defparam \Mux39~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N10
cycloneive_lcell_comb \Mux39~13 (
// Equation(s):
// \Mux39~13_combout  = (\prif.imemload_id [17] & ((\Mux39~12_combout  & ((\reg_file[7][24]~q ))) # (!\Mux39~12_combout  & (\reg_file[6][24]~q )))) # (!\prif.imemload_id [17] & (((\Mux39~12_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][24]~q ),
	.datac(\reg_file[7][24]~q ),
	.datad(\Mux39~12_combout ),
	.cin(gnd),
	.combout(\Mux39~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~13 .lut_mask = 16'hF588;
defparam \Mux39~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N15
dffeas \reg_file[1][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][24] .is_wysiwyg = "true";
defparam \reg_file[1][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N28
cycloneive_lcell_comb \reg_file[3][24]~feeder (
// Equation(s):
// \reg_file[3][24]~feeder_combout  = \reg_file_nxt[31][24]~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][24]~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[3][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[3][24]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[3][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N29
dffeas \reg_file[3][24] (
	.clk(!CLK),
	.d(\reg_file[3][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][24] .is_wysiwyg = "true";
defparam \reg_file[3][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N14
cycloneive_lcell_comb \Mux39~14 (
// Equation(s):
// \Mux39~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][24]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][24]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][24]~q ),
	.datad(\reg_file[3][24]~q ),
	.cin(gnd),
	.combout(\Mux39~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~14 .lut_mask = 16'hC840;
defparam \Mux39~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N29
dffeas \reg_file[2][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][24] .is_wysiwyg = "true";
defparam \reg_file[2][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N20
cycloneive_lcell_comb \Mux39~15 (
// Equation(s):
// \Mux39~15_combout  = (\Mux39~14_combout ) # ((\prif.imemload_id [17] & (!\prif.imemload_id [16] & \reg_file[2][24]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux39~14_combout ),
	.datad(\reg_file[2][24]~q ),
	.cin(gnd),
	.combout(\Mux39~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~15 .lut_mask = 16'hF2F0;
defparam \Mux39~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N30
cycloneive_lcell_comb \Mux39~16 (
// Equation(s):
// \Mux39~16_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\Mux39~13_combout )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\Mux39~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux39~13_combout ),
	.datad(\Mux39~15_combout ),
	.cin(gnd),
	.combout(\Mux39~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~16 .lut_mask = 16'hB9A8;
defparam \Mux39~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N11
dffeas \reg_file[11][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][24] .is_wysiwyg = "true";
defparam \reg_file[11][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N17
dffeas \reg_file[9][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][24] .is_wysiwyg = "true";
defparam \reg_file[9][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N11
dffeas \reg_file[8][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][24] .is_wysiwyg = "true";
defparam \reg_file[8][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N9
dffeas \reg_file[10][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][24] .is_wysiwyg = "true";
defparam \reg_file[10][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N10
cycloneive_lcell_comb \Mux39~10 (
// Equation(s):
// \Mux39~10_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][24]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][24]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[8][24]~q ),
	.datad(\reg_file[10][24]~q ),
	.cin(gnd),
	.combout(\Mux39~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~10 .lut_mask = 16'hDC98;
defparam \Mux39~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N16
cycloneive_lcell_comb \Mux39~11 (
// Equation(s):
// \Mux39~11_combout  = (\prif.imemload_id [16] & ((\Mux39~10_combout  & (\reg_file[11][24]~q )) # (!\Mux39~10_combout  & ((\reg_file[9][24]~q ))))) # (!\prif.imemload_id [16] & (((\Mux39~10_combout ))))

	.dataa(\reg_file[11][24]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[9][24]~q ),
	.datad(\Mux39~10_combout ),
	.cin(gnd),
	.combout(\Mux39~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~11 .lut_mask = 16'hBBC0;
defparam \Mux39~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N9
dffeas \reg_file[15][24] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][24]~84_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][24] .is_wysiwyg = "true";
defparam \reg_file[15][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N16
cycloneive_lcell_comb \reg_file[14][24]~feeder (
// Equation(s):
// \reg_file[14][24]~feeder_combout  = \reg_file_nxt[31][24]~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][24]~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[14][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][24]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[14][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N17
dffeas \reg_file[14][24] (
	.clk(!CLK),
	.d(\reg_file[14][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][24] .is_wysiwyg = "true";
defparam \reg_file[14][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N15
dffeas \reg_file[12][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][24] .is_wysiwyg = "true";
defparam \reg_file[12][24] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N29
dffeas \reg_file[13][24] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][24]~84_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][24] .is_wysiwyg = "true";
defparam \reg_file[13][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N28
cycloneive_lcell_comb \Mux39~17 (
// Equation(s):
// \Mux39~17_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][24]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][24]~q ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[12][24]~q ),
	.datac(\reg_file[13][24]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux39~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~17 .lut_mask = 16'hFA44;
defparam \Mux39~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N0
cycloneive_lcell_comb \Mux39~18 (
// Equation(s):
// \Mux39~18_combout  = (\prif.imemload_id [17] & ((\Mux39~17_combout  & (\reg_file[15][24]~q )) # (!\Mux39~17_combout  & ((\reg_file[14][24]~q ))))) # (!\prif.imemload_id [17] & (((\Mux39~17_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[15][24]~q ),
	.datac(\reg_file[14][24]~q ),
	.datad(\Mux39~17_combout ),
	.cin(gnd),
	.combout(\Mux39~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux39~18 .lut_mask = 16'hDDA0;
defparam \Mux39~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N2
cycloneive_lcell_comb \reg_file_nxt[31][16]~85 (
// Equation(s):
// \reg_file_nxt[31][16]~85_combout  = (\Mux148~1_combout  & (((\prif.regwrite_wb [2]) # (\prif.regwrite_wb [0])) # (!Equal8)))

	.dataa(Equal8),
	.datab(prifregwrite_wb_2),
	.datac(Mux148),
	.datad(prifregwrite_wb_0),
	.cin(gnd),
	.combout(\reg_file_nxt[31][16]~85_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][16]~85 .lut_mask = 16'hF0D0;
defparam \reg_file_nxt[31][16]~85 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N23
dffeas \reg_file[25][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][16] .is_wysiwyg = "true";
defparam \reg_file[25][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N14
cycloneive_lcell_comb \reg_file[29][16]~feeder (
// Equation(s):
// \reg_file[29][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][16]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][16]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N15
dffeas \reg_file[29][16] (
	.clk(!CLK),
	.d(\reg_file[29][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][16] .is_wysiwyg = "true";
defparam \reg_file[29][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N5
dffeas \reg_file[17][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][16] .is_wysiwyg = "true";
defparam \reg_file[17][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N4
cycloneive_lcell_comb \Mux47~0 (
// Equation(s):
// \Mux47~0_combout  = (\prif.imemload_id [18] & ((\reg_file[21][16]~q ) # ((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (((\reg_file[17][16]~q  & !\prif.imemload_id [19]))))

	.dataa(\reg_file[21][16]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[17][16]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux47~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~0 .lut_mask = 16'hCCB8;
defparam \Mux47~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N20
cycloneive_lcell_comb \Mux47~1 (
// Equation(s):
// \Mux47~1_combout  = (\prif.imemload_id [19] & ((\Mux47~0_combout  & ((\reg_file[29][16]~q ))) # (!\Mux47~0_combout  & (\reg_file[25][16]~q )))) # (!\prif.imemload_id [19] & (((\Mux47~0_combout ))))

	.dataa(\reg_file[25][16]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[29][16]~q ),
	.datad(\Mux47~0_combout ),
	.cin(gnd),
	.combout(\Mux47~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~1 .lut_mask = 16'hF388;
defparam \Mux47~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N6
cycloneive_lcell_comb \reg_file[31][16]~feeder (
// Equation(s):
// \reg_file[31][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][16]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[31][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][16]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[31][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N7
dffeas \reg_file[31][16] (
	.clk(!CLK),
	.d(\reg_file[31][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][16] .is_wysiwyg = "true";
defparam \reg_file[31][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N22
cycloneive_lcell_comb \reg_file[27][16]~feeder (
// Equation(s):
// \reg_file[27][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][16]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[27][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[27][16]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[27][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N23
dffeas \reg_file[27][16] (
	.clk(!CLK),
	.d(\reg_file[27][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][16] .is_wysiwyg = "true";
defparam \reg_file[27][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y26_N17
dffeas \reg_file[23][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][16] .is_wysiwyg = "true";
defparam \reg_file[23][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N16
cycloneive_lcell_comb \Mux47~7 (
// Equation(s):
// \Mux47~7_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[23][16]~q ))) # (!\prif.imemload_id [18] & (\reg_file[19][16]~q ))))

	.dataa(\reg_file[19][16]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][16]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux47~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~7 .lut_mask = 16'hFC22;
defparam \Mux47~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N12
cycloneive_lcell_comb \Mux47~8 (
// Equation(s):
// \Mux47~8_combout  = (\prif.imemload_id [19] & ((\Mux47~7_combout  & (\reg_file[31][16]~q )) # (!\Mux47~7_combout  & ((\reg_file[27][16]~q ))))) # (!\prif.imemload_id [19] & (((\Mux47~7_combout ))))

	.dataa(\reg_file[31][16]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][16]~q ),
	.datad(\Mux47~7_combout ),
	.cin(gnd),
	.combout(\Mux47~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~8 .lut_mask = 16'hBBC0;
defparam \Mux47~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N19
dffeas \reg_file[28][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][16] .is_wysiwyg = "true";
defparam \reg_file[28][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N21
dffeas \reg_file[20][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][16] .is_wysiwyg = "true";
defparam \reg_file[20][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N12
cycloneive_lcell_comb \reg_file[24][16]~feeder (
// Equation(s):
// \reg_file[24][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][16]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[24][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][16]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[24][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N13
dffeas \reg_file[24][16] (
	.clk(!CLK),
	.d(\reg_file[24][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][16] .is_wysiwyg = "true";
defparam \reg_file[24][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N27
dffeas \reg_file[16][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][16] .is_wysiwyg = "true";
defparam \reg_file[16][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N26
cycloneive_lcell_comb \Mux47~4 (
// Equation(s):
// \Mux47~4_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[24][16]~q )) # (!\prif.imemload_id [19] & ((\reg_file[16][16]~q )))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[24][16]~q ),
	.datac(\reg_file[16][16]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux47~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~4 .lut_mask = 16'hEE50;
defparam \Mux47~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N14
cycloneive_lcell_comb \Mux47~5 (
// Equation(s):
// \Mux47~5_combout  = (\prif.imemload_id [18] & ((\Mux47~4_combout  & (\reg_file[28][16]~q )) # (!\Mux47~4_combout  & ((\reg_file[20][16]~q ))))) # (!\prif.imemload_id [18] & (((\Mux47~4_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[28][16]~q ),
	.datac(\reg_file[20][16]~q ),
	.datad(\Mux47~4_combout ),
	.cin(gnd),
	.combout(\Mux47~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~5 .lut_mask = 16'hDDA0;
defparam \Mux47~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N3
dffeas \reg_file[30][16] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][16]~85_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][16] .is_wysiwyg = "true";
defparam \reg_file[30][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N8
cycloneive_lcell_comb \reg_file[22][16]~feeder (
// Equation(s):
// \reg_file[22][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][16]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[22][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][16]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[22][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N9
dffeas \reg_file[22][16] (
	.clk(!CLK),
	.d(\reg_file[22][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][16] .is_wysiwyg = "true";
defparam \reg_file[22][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N28
cycloneive_lcell_comb \Mux47~3 (
// Equation(s):
// \Mux47~3_combout  = (\Mux47~2_combout  & ((\reg_file[30][16]~q ) # ((!\prif.imemload_id [18])))) # (!\Mux47~2_combout  & (((\reg_file[22][16]~q  & \prif.imemload_id [18]))))

	.dataa(\Mux47~2_combout ),
	.datab(\reg_file[30][16]~q ),
	.datac(\reg_file[22][16]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux47~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~3 .lut_mask = 16'hD8AA;
defparam \Mux47~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y31_N20
cycloneive_lcell_comb \Mux47~6 (
// Equation(s):
// \Mux47~6_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16]) # (\Mux47~3_combout )))) # (!\prif.imemload_id [17] & (\Mux47~5_combout  & (!\prif.imemload_id [16])))

	.dataa(prifimemload_id_17),
	.datab(\Mux47~5_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux47~3_combout ),
	.cin(gnd),
	.combout(\Mux47~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~6 .lut_mask = 16'hAEA4;
defparam \Mux47~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N29
dffeas \reg_file[1][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][16] .is_wysiwyg = "true";
defparam \reg_file[1][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N28
cycloneive_lcell_comb \Mux47~14 (
// Equation(s):
// \Mux47~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][16]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][16]~q )))))

	.dataa(\reg_file[3][16]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[1][16]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux47~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~14 .lut_mask = 16'hB800;
defparam \Mux47~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y27_N7
dffeas \reg_file[2][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][16] .is_wysiwyg = "true";
defparam \reg_file[2][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N14
cycloneive_lcell_comb \Mux47~15 (
// Equation(s):
// \Mux47~15_combout  = (\Mux47~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][16]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\Mux47~14_combout ),
	.datad(\reg_file[2][16]~q ),
	.cin(gnd),
	.combout(\Mux47~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~15 .lut_mask = 16'hF4F0;
defparam \Mux47~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N9
dffeas \reg_file[6][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][16] .is_wysiwyg = "true";
defparam \reg_file[6][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N19
dffeas \reg_file[7][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][16] .is_wysiwyg = "true";
defparam \reg_file[7][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N19
dffeas \reg_file[4][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][16] .is_wysiwyg = "true";
defparam \reg_file[4][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N29
dffeas \reg_file[5][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][16] .is_wysiwyg = "true";
defparam \reg_file[5][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N18
cycloneive_lcell_comb \Mux47~12 (
// Equation(s):
// \Mux47~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][16]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][16]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][16]~q ),
	.datad(\reg_file[5][16]~q ),
	.cin(gnd),
	.combout(\Mux47~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~12 .lut_mask = 16'hBA98;
defparam \Mux47~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N18
cycloneive_lcell_comb \Mux47~13 (
// Equation(s):
// \Mux47~13_combout  = (\prif.imemload_id [17] & ((\Mux47~12_combout  & ((\reg_file[7][16]~q ))) # (!\Mux47~12_combout  & (\reg_file[6][16]~q )))) # (!\prif.imemload_id [17] & (((\Mux47~12_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][16]~q ),
	.datac(\reg_file[7][16]~q ),
	.datad(\Mux47~12_combout ),
	.cin(gnd),
	.combout(\Mux47~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~13 .lut_mask = 16'hF588;
defparam \Mux47~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N20
cycloneive_lcell_comb \Mux47~16 (
// Equation(s):
// \Mux47~16_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\Mux47~13_combout ))) # (!\prif.imemload_id [18] & (\Mux47~15_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\Mux47~15_combout ),
	.datac(prifimemload_id_18),
	.datad(\Mux47~13_combout ),
	.cin(gnd),
	.combout(\Mux47~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~16 .lut_mask = 16'hF4A4;
defparam \Mux47~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N15
dffeas \reg_file[12][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][16] .is_wysiwyg = "true";
defparam \reg_file[12][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N25
dffeas \reg_file[13][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][16] .is_wysiwyg = "true";
defparam \reg_file[13][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N14
cycloneive_lcell_comb \Mux47~17 (
// Equation(s):
// \Mux47~17_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[13][16]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[12][16]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[12][16]~q ),
	.datad(\reg_file[13][16]~q ),
	.cin(gnd),
	.combout(\Mux47~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~17 .lut_mask = 16'hBA98;
defparam \Mux47~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N1
dffeas \reg_file[14][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][16] .is_wysiwyg = "true";
defparam \reg_file[14][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N24
cycloneive_lcell_comb \reg_file[15][16]~feeder (
// Equation(s):
// \reg_file[15][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][16]~85_combout ),
	.cin(gnd),
	.combout(\reg_file[15][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[15][16]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[15][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N25
dffeas \reg_file[15][16] (
	.clk(!CLK),
	.d(\reg_file[15][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][16] .is_wysiwyg = "true";
defparam \reg_file[15][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N26
cycloneive_lcell_comb \Mux47~18 (
// Equation(s):
// \Mux47~18_combout  = (\Mux47~17_combout  & (((\reg_file[15][16]~q ) # (!\prif.imemload_id [17])))) # (!\Mux47~17_combout  & (\reg_file[14][16]~q  & (\prif.imemload_id [17])))

	.dataa(\Mux47~17_combout ),
	.datab(\reg_file[14][16]~q ),
	.datac(prifimemload_id_17),
	.datad(\reg_file[15][16]~q ),
	.cin(gnd),
	.combout(\Mux47~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~18 .lut_mask = 16'hEA4A;
defparam \Mux47~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N6
cycloneive_lcell_comb \reg_file[9][16]~feeder (
// Equation(s):
// \reg_file[9][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][16]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[9][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[9][16]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[9][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N7
dffeas \reg_file[9][16] (
	.clk(!CLK),
	.d(\reg_file[9][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][16] .is_wysiwyg = "true";
defparam \reg_file[9][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N19
dffeas \reg_file[8][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][16] .is_wysiwyg = "true";
defparam \reg_file[8][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N21
dffeas \reg_file[10][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][16] .is_wysiwyg = "true";
defparam \reg_file[10][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N20
cycloneive_lcell_comb \Mux47~10 (
// Equation(s):
// \Mux47~10_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][16]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][16]~q ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[8][16]~q ),
	.datac(\reg_file[10][16]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux47~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~10 .lut_mask = 16'hFA44;
defparam \Mux47~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N8
cycloneive_lcell_comb \reg_file[11][16]~feeder (
// Equation(s):
// \reg_file[11][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][16]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[11][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[11][16]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[11][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y27_N9
dffeas \reg_file[11][16] (
	.clk(!CLK),
	.d(\reg_file[11][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][16] .is_wysiwyg = "true";
defparam \reg_file[11][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N8
cycloneive_lcell_comb \Mux47~11 (
// Equation(s):
// \Mux47~11_combout  = (\Mux47~10_combout  & (((\reg_file[11][16]~q ) # (!\prif.imemload_id [16])))) # (!\Mux47~10_combout  & (\reg_file[9][16]~q  & ((\prif.imemload_id [16]))))

	.dataa(\reg_file[9][16]~q ),
	.datab(\Mux47~10_combout ),
	.datac(\reg_file[11][16]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux47~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux47~11 .lut_mask = 16'hE2CC;
defparam \Mux47~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N0
cycloneive_lcell_comb \reg_file_nxt[31][19]~86 (
// Equation(s):
// \reg_file_nxt[31][19]~86_combout  = (\Mux145~1_combout  & ((\prif.regwrite_wb [0]) # ((\prif.regwrite_wb [2]) # (!Equal8))))

	.dataa(Mux145),
	.datab(prifregwrite_wb_0),
	.datac(Equal8),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\reg_file_nxt[31][19]~86_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][19]~86 .lut_mask = 16'hAA8A;
defparam \reg_file_nxt[31][19]~86 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N20
cycloneive_lcell_comb \reg_file[29][19]~feeder (
// Equation(s):
// \reg_file[29][19]~feeder_combout  = \reg_file_nxt[31][19]~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][19]~86_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][19]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N21
dffeas \reg_file[29][19] (
	.clk(!CLK),
	.d(\reg_file[29][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][19] .is_wysiwyg = "true";
defparam \reg_file[29][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N4
cycloneive_lcell_comb \reg_file[21][19]~feeder (
// Equation(s):
// \reg_file[21][19]~feeder_combout  = \reg_file_nxt[31][19]~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][19]~86_combout ),
	.cin(gnd),
	.combout(\reg_file[21][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][19]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[21][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N5
dffeas \reg_file[21][19] (
	.clk(!CLK),
	.d(\reg_file[21][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][19] .is_wysiwyg = "true";
defparam \reg_file[21][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N27
dffeas \reg_file[17][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][19] .is_wysiwyg = "true";
defparam \reg_file[17][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y28_N17
dffeas \reg_file[25][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][19] .is_wysiwyg = "true";
defparam \reg_file[25][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N26
cycloneive_lcell_comb \Mux44~0 (
// Equation(s):
// \Mux44~0_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[25][19]~q ))) # (!\prif.imemload_id [19] & (\reg_file[17][19]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][19]~q ),
	.datad(\reg_file[25][19]~q ),
	.cin(gnd),
	.combout(\Mux44~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~0 .lut_mask = 16'hDC98;
defparam \Mux44~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N18
cycloneive_lcell_comb \Mux44~1 (
// Equation(s):
// \Mux44~1_combout  = (\prif.imemload_id [18] & ((\Mux44~0_combout  & (\reg_file[29][19]~q )) # (!\Mux44~0_combout  & ((\reg_file[21][19]~q ))))) # (!\prif.imemload_id [18] & (((\Mux44~0_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[29][19]~q ),
	.datac(\reg_file[21][19]~q ),
	.datad(\Mux44~0_combout ),
	.cin(gnd),
	.combout(\Mux44~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~1 .lut_mask = 16'hDDA0;
defparam \Mux44~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N4
cycloneive_lcell_comb \reg_file[20][19]~feeder (
// Equation(s):
// \reg_file[20][19]~feeder_combout  = \reg_file_nxt[31][19]~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][19]~86_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[20][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[20][19]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[20][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N5
dffeas \reg_file[20][19] (
	.clk(!CLK),
	.d(\reg_file[20][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][19] .is_wysiwyg = "true";
defparam \reg_file[20][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N15
dffeas \reg_file[16][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][19] .is_wysiwyg = "true";
defparam \reg_file[16][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N14
cycloneive_lcell_comb \Mux44~4 (
// Equation(s):
// \Mux44~4_combout  = (\prif.imemload_id [18] & ((\reg_file[20][19]~q ) # ((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (((\reg_file[16][19]~q  & !\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[20][19]~q ),
	.datac(\reg_file[16][19]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux44~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~4 .lut_mask = 16'hAAD8;
defparam \Mux44~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N11
dffeas \reg_file[28][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][19] .is_wysiwyg = "true";
defparam \reg_file[28][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N8
cycloneive_lcell_comb \Mux44~5 (
// Equation(s):
// \Mux44~5_combout  = (\Mux44~4_combout  & (((\reg_file[28][19]~q ) # (!\prif.imemload_id [19])))) # (!\Mux44~4_combout  & (\reg_file[24][19]~q  & (\prif.imemload_id [19])))

	.dataa(\reg_file[24][19]~q ),
	.datab(\Mux44~4_combout ),
	.datac(prifimemload_id_19),
	.datad(\reg_file[28][19]~q ),
	.cin(gnd),
	.combout(\Mux44~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~5 .lut_mask = 16'hEC2C;
defparam \Mux44~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N23
dffeas \reg_file[22][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][19] .is_wysiwyg = "true";
defparam \reg_file[22][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N23
dffeas \reg_file[18][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][19] .is_wysiwyg = "true";
defparam \reg_file[18][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N22
cycloneive_lcell_comb \Mux44~2 (
// Equation(s):
// \Mux44~2_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[22][19]~q )) # (!\prif.imemload_id [18] & ((\reg_file[18][19]~q )))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[22][19]~q ),
	.datad(\reg_file[18][19]~q ),
	.cin(gnd),
	.combout(\Mux44~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~2 .lut_mask = 16'hD9C8;
defparam \Mux44~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N23
dffeas \reg_file[30][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][19] .is_wysiwyg = "true";
defparam \reg_file[30][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N22
cycloneive_lcell_comb \Mux44~3 (
// Equation(s):
// \Mux44~3_combout  = (\Mux44~2_combout  & (((\reg_file[30][19]~q ) # (!\prif.imemload_id [19])))) # (!\Mux44~2_combout  & (\reg_file[26][19]~q  & ((\prif.imemload_id [19]))))

	.dataa(\reg_file[26][19]~q ),
	.datab(\Mux44~2_combout ),
	.datac(\reg_file[30][19]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux44~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~3 .lut_mask = 16'hE2CC;
defparam \Mux44~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N14
cycloneive_lcell_comb \Mux44~6 (
// Equation(s):
// \Mux44~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux44~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & (\Mux44~5_combout )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux44~5_combout ),
	.datad(\Mux44~3_combout ),
	.cin(gnd),
	.combout(\Mux44~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~6 .lut_mask = 16'hBA98;
defparam \Mux44~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N15
dffeas \reg_file[19][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][19] .is_wysiwyg = "true";
defparam \reg_file[19][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N1
dffeas \reg_file[27][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][19] .is_wysiwyg = "true";
defparam \reg_file[27][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N0
cycloneive_lcell_comb \Mux44~7 (
// Equation(s):
// \Mux44~7_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[27][19]~q ))) # (!\prif.imemload_id [19] & (\reg_file[19][19]~q ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[19][19]~q ),
	.datac(\reg_file[27][19]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux44~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~7 .lut_mask = 16'hFA44;
defparam \Mux44~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N26
cycloneive_lcell_comb \reg_file[23][19]~feeder (
// Equation(s):
// \reg_file[23][19]~feeder_combout  = \reg_file_nxt[31][19]~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][19]~86_combout ),
	.cin(gnd),
	.combout(\reg_file[23][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][19]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[23][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N27
dffeas \reg_file[23][19] (
	.clk(!CLK),
	.d(\reg_file[23][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][19] .is_wysiwyg = "true";
defparam \reg_file[23][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N28
cycloneive_lcell_comb \reg_file[31][19]~feeder (
// Equation(s):
// \reg_file[31][19]~feeder_combout  = \reg_file_nxt[31][19]~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][19]~86_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[31][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][19]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[31][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y32_N29
dffeas \reg_file[31][19] (
	.clk(!CLK),
	.d(\reg_file[31][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][19] .is_wysiwyg = "true";
defparam \reg_file[31][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N18
cycloneive_lcell_comb \Mux44~8 (
// Equation(s):
// \Mux44~8_combout  = (\Mux44~7_combout  & (((\reg_file[31][19]~q ) # (!\prif.imemload_id [18])))) # (!\Mux44~7_combout  & (\reg_file[23][19]~q  & (\prif.imemload_id [18])))

	.dataa(\Mux44~7_combout ),
	.datab(\reg_file[23][19]~q ),
	.datac(prifimemload_id_18),
	.datad(\reg_file[31][19]~q ),
	.cin(gnd),
	.combout(\Mux44~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~8 .lut_mask = 16'hEA4A;
defparam \Mux44~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N26
cycloneive_lcell_comb \reg_file[6][19]~feeder (
// Equation(s):
// \reg_file[6][19]~feeder_combout  = \reg_file_nxt[31][19]~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][19]~86_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][19]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N27
dffeas \reg_file[6][19] (
	.clk(!CLK),
	.d(\reg_file[6][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][19] .is_wysiwyg = "true";
defparam \reg_file[6][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N1
dffeas \reg_file[7][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][19] .is_wysiwyg = "true";
defparam \reg_file[7][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N11
dffeas \reg_file[4][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][19] .is_wysiwyg = "true";
defparam \reg_file[4][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N1
dffeas \reg_file[5][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][19] .is_wysiwyg = "true";
defparam \reg_file[5][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N10
cycloneive_lcell_comb \Mux44~10 (
// Equation(s):
// \Mux44~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][19]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][19]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][19]~q ),
	.datad(\reg_file[5][19]~q ),
	.cin(gnd),
	.combout(\Mux44~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~10 .lut_mask = 16'hBA98;
defparam \Mux44~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N0
cycloneive_lcell_comb \Mux44~11 (
// Equation(s):
// \Mux44~11_combout  = (\prif.imemload_id [17] & ((\Mux44~10_combout  & ((\reg_file[7][19]~q ))) # (!\Mux44~10_combout  & (\reg_file[6][19]~q )))) # (!\prif.imemload_id [17] & (((\Mux44~10_combout ))))

	.dataa(\reg_file[6][19]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[7][19]~q ),
	.datad(\Mux44~10_combout ),
	.cin(gnd),
	.combout(\Mux44~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~11 .lut_mask = 16'hF388;
defparam \Mux44~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N1
dffeas \reg_file[15][19] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][19]~86_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][19] .is_wysiwyg = "true";
defparam \reg_file[15][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N3
dffeas \reg_file[12][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][19] .is_wysiwyg = "true";
defparam \reg_file[12][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N21
dffeas \reg_file[13][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][19] .is_wysiwyg = "true";
defparam \reg_file[13][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N2
cycloneive_lcell_comb \Mux44~17 (
// Equation(s):
// \Mux44~17_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[13][19]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[12][19]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[12][19]~q ),
	.datad(\reg_file[13][19]~q ),
	.cin(gnd),
	.combout(\Mux44~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~17 .lut_mask = 16'hBA98;
defparam \Mux44~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y26_N19
dffeas \reg_file[14][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][19] .is_wysiwyg = "true";
defparam \reg_file[14][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N30
cycloneive_lcell_comb \Mux44~18 (
// Equation(s):
// \Mux44~18_combout  = (\prif.imemload_id [17] & ((\Mux44~17_combout  & (\reg_file[15][19]~q )) # (!\Mux44~17_combout  & ((\reg_file[14][19]~q ))))) # (!\prif.imemload_id [17] & (((\Mux44~17_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[15][19]~q ),
	.datac(\Mux44~17_combout ),
	.datad(\reg_file[14][19]~q ),
	.cin(gnd),
	.combout(\Mux44~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~18 .lut_mask = 16'hDAD0;
defparam \Mux44~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N3
dffeas \reg_file[3][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][19] .is_wysiwyg = "true";
defparam \reg_file[3][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N9
dffeas \reg_file[1][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][19] .is_wysiwyg = "true";
defparam \reg_file[1][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N8
cycloneive_lcell_comb \Mux44~14 (
// Equation(s):
// \Mux44~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][19]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][19]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[3][19]~q ),
	.datac(\reg_file[1][19]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux44~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~14 .lut_mask = 16'hD800;
defparam \Mux44~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N20
cycloneive_lcell_comb \reg_file[2][19]~feeder (
// Equation(s):
// \reg_file[2][19]~feeder_combout  = \reg_file_nxt[31][19]~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][19]~86_combout ),
	.cin(gnd),
	.combout(\reg_file[2][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][19]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[2][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N21
dffeas \reg_file[2][19] (
	.clk(!CLK),
	.d(\reg_file[2][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][19] .is_wysiwyg = "true";
defparam \reg_file[2][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N6
cycloneive_lcell_comb \Mux44~15 (
// Equation(s):
// \Mux44~15_combout  = (\Mux44~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][19]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\Mux44~14_combout ),
	.datad(\reg_file[2][19]~q ),
	.cin(gnd),
	.combout(\Mux44~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~15 .lut_mask = 16'hF4F0;
defparam \Mux44~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N25
dffeas \reg_file[10][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][19] .is_wysiwyg = "true";
defparam \reg_file[10][19] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N27
dffeas \reg_file[8][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][19] .is_wysiwyg = "true";
defparam \reg_file[8][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N26
cycloneive_lcell_comb \Mux44~12 (
// Equation(s):
// \Mux44~12_combout  = (\prif.imemload_id [17] & ((\reg_file[10][19]~q ) # ((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (((\reg_file[8][19]~q  & !\prif.imemload_id [16]))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[10][19]~q ),
	.datac(\reg_file[8][19]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux44~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~12 .lut_mask = 16'hAAD8;
defparam \Mux44~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N5
dffeas \reg_file[9][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][19] .is_wysiwyg = "true";
defparam \reg_file[9][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N22
cycloneive_lcell_comb \Mux44~13 (
// Equation(s):
// \Mux44~13_combout  = (\Mux44~12_combout  & ((\reg_file[11][19]~q ) # ((!\prif.imemload_id [16])))) # (!\Mux44~12_combout  & (((\reg_file[9][19]~q  & \prif.imemload_id [16]))))

	.dataa(\reg_file[11][19]~q ),
	.datab(\Mux44~12_combout ),
	.datac(\reg_file[9][19]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux44~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~13 .lut_mask = 16'hB8CC;
defparam \Mux44~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N28
cycloneive_lcell_comb \Mux44~16 (
// Equation(s):
// \Mux44~16_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\Mux44~13_combout ))) # (!\prif.imemload_id [19] & (\Mux44~15_combout ))))

	.dataa(\Mux44~15_combout ),
	.datab(prifimemload_id_18),
	.datac(\Mux44~13_combout ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux44~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux44~16 .lut_mask = 16'hFC22;
defparam \Mux44~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N8
cycloneive_lcell_comb \reg_file_nxt[31][17]~87 (
// Equation(s):
// \reg_file_nxt[31][17]~87_combout  = (\Mux147~1_combout  & (((\prif.regwrite_wb [2]) # (\prif.regwrite_wb [0])) # (!Equal8)))

	.dataa(Equal8),
	.datab(prifregwrite_wb_2),
	.datac(Mux147),
	.datad(prifregwrite_wb_0),
	.cin(gnd),
	.combout(\reg_file_nxt[31][17]~87_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][17]~87 .lut_mask = 16'hF0D0;
defparam \reg_file_nxt[31][17]~87 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N11
dffeas \reg_file[29][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][17] .is_wysiwyg = "true";
defparam \reg_file[29][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N21
dffeas \reg_file[17][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][17] .is_wysiwyg = "true";
defparam \reg_file[17][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N4
cycloneive_lcell_comb \reg_file[25][17]~feeder (
// Equation(s):
// \reg_file[25][17]~feeder_combout  = \reg_file_nxt[31][17]~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][17]~87_combout ),
	.cin(gnd),
	.combout(\reg_file[25][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][17]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[25][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N5
dffeas \reg_file[25][17] (
	.clk(!CLK),
	.d(\reg_file[25][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][17] .is_wysiwyg = "true";
defparam \reg_file[25][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N20
cycloneive_lcell_comb \Mux46~0 (
// Equation(s):
// \Mux46~0_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[25][17]~q ))) # (!\prif.imemload_id [19] & (\reg_file[17][17]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][17]~q ),
	.datad(\reg_file[25][17]~q ),
	.cin(gnd),
	.combout(\Mux46~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~0 .lut_mask = 16'hDC98;
defparam \Mux46~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N22
cycloneive_lcell_comb \reg_file[21][17]~feeder (
// Equation(s):
// \reg_file[21][17]~feeder_combout  = \reg_file_nxt[31][17]~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][17]~87_combout ),
	.cin(gnd),
	.combout(\reg_file[21][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][17]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[21][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N23
dffeas \reg_file[21][17] (
	.clk(!CLK),
	.d(\reg_file[21][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][17] .is_wysiwyg = "true";
defparam \reg_file[21][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N8
cycloneive_lcell_comb \Mux46~1 (
// Equation(s):
// \Mux46~1_combout  = (\prif.imemload_id [18] & ((\Mux46~0_combout  & (\reg_file[29][17]~q )) # (!\Mux46~0_combout  & ((\reg_file[21][17]~q ))))) # (!\prif.imemload_id [18] & (((\Mux46~0_combout ))))

	.dataa(\reg_file[29][17]~q ),
	.datab(prifimemload_id_18),
	.datac(\Mux46~0_combout ),
	.datad(\reg_file[21][17]~q ),
	.cin(gnd),
	.combout(\Mux46~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~1 .lut_mask = 16'hBCB0;
defparam \Mux46~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N12
cycloneive_lcell_comb \reg_file[23][17]~feeder (
// Equation(s):
// \reg_file[23][17]~feeder_combout  = \reg_file_nxt[31][17]~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][17]~87_combout ),
	.cin(gnd),
	.combout(\reg_file[23][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][17]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[23][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N13
dffeas \reg_file[23][17] (
	.clk(!CLK),
	.d(\reg_file[23][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][17] .is_wysiwyg = "true";
defparam \reg_file[23][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N23
dffeas \reg_file[31][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][17] .is_wysiwyg = "true";
defparam \reg_file[31][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N25
dffeas \reg_file[27][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][17] .is_wysiwyg = "true";
defparam \reg_file[27][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N3
dffeas \reg_file[19][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][17] .is_wysiwyg = "true";
defparam \reg_file[19][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N24
cycloneive_lcell_comb \Mux46~7 (
// Equation(s):
// \Mux46~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][17]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][17]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][17]~q ),
	.datad(\reg_file[19][17]~q ),
	.cin(gnd),
	.combout(\Mux46~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~7 .lut_mask = 16'hD9C8;
defparam \Mux46~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N22
cycloneive_lcell_comb \Mux46~8 (
// Equation(s):
// \Mux46~8_combout  = (\prif.imemload_id [18] & ((\Mux46~7_combout  & ((\reg_file[31][17]~q ))) # (!\Mux46~7_combout  & (\reg_file[23][17]~q )))) # (!\prif.imemload_id [18] & (((\Mux46~7_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[23][17]~q ),
	.datac(\reg_file[31][17]~q ),
	.datad(\Mux46~7_combout ),
	.cin(gnd),
	.combout(\Mux46~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~8 .lut_mask = 16'hF588;
defparam \Mux46~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N1
dffeas \reg_file[30][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][17] .is_wysiwyg = "true";
defparam \reg_file[30][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N1
dffeas \reg_file[22][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][17] .is_wysiwyg = "true";
defparam \reg_file[22][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N7
dffeas \reg_file[18][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][17] .is_wysiwyg = "true";
defparam \reg_file[18][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N0
cycloneive_lcell_comb \Mux46~2 (
// Equation(s):
// \Mux46~2_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[22][17]~q )) # (!\prif.imemload_id [18] & ((\reg_file[18][17]~q )))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[22][17]~q ),
	.datad(\reg_file[18][17]~q ),
	.cin(gnd),
	.combout(\Mux46~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~2 .lut_mask = 16'hD9C8;
defparam \Mux46~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N0
cycloneive_lcell_comb \Mux46~3 (
// Equation(s):
// \Mux46~3_combout  = (\prif.imemload_id [19] & ((\Mux46~2_combout  & ((\reg_file[30][17]~q ))) # (!\Mux46~2_combout  & (\reg_file[26][17]~q )))) # (!\prif.imemload_id [19] & (((\Mux46~2_combout ))))

	.dataa(\reg_file[26][17]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[30][17]~q ),
	.datad(\Mux46~2_combout ),
	.cin(gnd),
	.combout(\Mux46~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~3 .lut_mask = 16'hF388;
defparam \Mux46~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N17
dffeas \reg_file[24][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][17] .is_wysiwyg = "true";
defparam \reg_file[24][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N27
dffeas \reg_file[28][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][17] .is_wysiwyg = "true";
defparam \reg_file[28][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N16
cycloneive_lcell_comb \Mux46~5 (
// Equation(s):
// \Mux46~5_combout  = (\Mux46~4_combout  & (((\reg_file[28][17]~q )) # (!\prif.imemload_id [19]))) # (!\Mux46~4_combout  & (\prif.imemload_id [19] & (\reg_file[24][17]~q )))

	.dataa(\Mux46~4_combout ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[24][17]~q ),
	.datad(\reg_file[28][17]~q ),
	.cin(gnd),
	.combout(\Mux46~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~5 .lut_mask = 16'hEA62;
defparam \Mux46~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N18
cycloneive_lcell_comb \Mux46~6 (
// Equation(s):
// \Mux46~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux46~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & ((\Mux46~5_combout ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux46~3_combout ),
	.datad(\Mux46~5_combout ),
	.cin(gnd),
	.combout(\Mux46~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~6 .lut_mask = 16'hB9A8;
defparam \Mux46~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N30
cycloneive_lcell_comb \reg_file[9][17]~feeder (
// Equation(s):
// \reg_file[9][17]~feeder_combout  = \reg_file_nxt[31][17]~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][17]~87_combout ),
	.cin(gnd),
	.combout(\reg_file[9][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[9][17]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[9][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N31
dffeas \reg_file[9][17] (
	.clk(!CLK),
	.d(\reg_file[9][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][17] .is_wysiwyg = "true";
defparam \reg_file[9][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N21
dffeas \reg_file[10][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][17] .is_wysiwyg = "true";
defparam \reg_file[10][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N23
dffeas \reg_file[8][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][17] .is_wysiwyg = "true";
defparam \reg_file[8][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N22
cycloneive_lcell_comb \Mux46~12 (
// Equation(s):
// \Mux46~12_combout  = (\prif.imemload_id [17] & ((\reg_file[10][17]~q ) # ((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (((\reg_file[8][17]~q  & !\prif.imemload_id [16]))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[10][17]~q ),
	.datac(\reg_file[8][17]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux46~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~12 .lut_mask = 16'hAAD8;
defparam \Mux46~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N4
cycloneive_lcell_comb \Mux46~13 (
// Equation(s):
// \Mux46~13_combout  = (\prif.imemload_id [16] & ((\Mux46~12_combout  & (\reg_file[11][17]~q )) # (!\Mux46~12_combout  & ((\reg_file[9][17]~q ))))) # (!\prif.imemload_id [16] & (((\Mux46~12_combout ))))

	.dataa(\reg_file[11][17]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[9][17]~q ),
	.datad(\Mux46~12_combout ),
	.cin(gnd),
	.combout(\Mux46~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~13 .lut_mask = 16'hBBC0;
defparam \Mux46~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N27
dffeas \reg_file[1][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][17] .is_wysiwyg = "true";
defparam \reg_file[1][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N24
cycloneive_lcell_comb \reg_file[3][17]~feeder (
// Equation(s):
// \reg_file[3][17]~feeder_combout  = \reg_file_nxt[31][17]~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][17]~87_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[3][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[3][17]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[3][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N25
dffeas \reg_file[3][17] (
	.clk(!CLK),
	.d(\reg_file[3][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][17] .is_wysiwyg = "true";
defparam \reg_file[3][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N16
cycloneive_lcell_comb \Mux46~14 (
// Equation(s):
// \Mux46~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][17]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][17]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][17]~q ),
	.datad(\reg_file[3][17]~q ),
	.cin(gnd),
	.combout(\Mux46~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~14 .lut_mask = 16'hC840;
defparam \Mux46~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N20
cycloneive_lcell_comb \Mux46~15 (
// Equation(s):
// \Mux46~15_combout  = (\Mux46~14_combout ) # ((\reg_file[2][17]~q  & (!\prif.imemload_id [16] & \prif.imemload_id [17])))

	.dataa(\reg_file[2][17]~q ),
	.datab(prifimemload_id_16),
	.datac(prifimemload_id_17),
	.datad(\Mux46~14_combout ),
	.cin(gnd),
	.combout(\Mux46~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~15 .lut_mask = 16'hFF20;
defparam \Mux46~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N10
cycloneive_lcell_comb \Mux46~16 (
// Equation(s):
// \Mux46~16_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\Mux46~13_combout )) # (!\prif.imemload_id [19] & ((\Mux46~15_combout )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux46~13_combout ),
	.datad(\Mux46~15_combout ),
	.cin(gnd),
	.combout(\Mux46~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~16 .lut_mask = 16'hD9C8;
defparam \Mux46~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N9
dffeas \reg_file[13][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][17] .is_wysiwyg = "true";
defparam \reg_file[13][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N7
dffeas \reg_file[12][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][17] .is_wysiwyg = "true";
defparam \reg_file[12][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N8
cycloneive_lcell_comb \Mux46~17 (
// Equation(s):
// \Mux46~17_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[13][17]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[12][17]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[13][17]~q ),
	.datad(\reg_file[12][17]~q ),
	.cin(gnd),
	.combout(\Mux46~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~17 .lut_mask = 16'hB9A8;
defparam \Mux46~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N29
dffeas \reg_file[14][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][17] .is_wysiwyg = "true";
defparam \reg_file[14][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N9
dffeas \reg_file[15][17] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][17]~87_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][17] .is_wysiwyg = "true";
defparam \reg_file[15][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N28
cycloneive_lcell_comb \Mux46~18 (
// Equation(s):
// \Mux46~18_combout  = (\Mux46~17_combout  & (((\reg_file[15][17]~q )) # (!\prif.imemload_id [17]))) # (!\Mux46~17_combout  & (\prif.imemload_id [17] & (\reg_file[14][17]~q )))

	.dataa(\Mux46~17_combout ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[14][17]~q ),
	.datad(\reg_file[15][17]~q ),
	.cin(gnd),
	.combout(\Mux46~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~18 .lut_mask = 16'hEA62;
defparam \Mux46~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y29_N23
dffeas \reg_file[7][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][17] .is_wysiwyg = "true";
defparam \reg_file[7][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y29_N1
dffeas \reg_file[6][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][17] .is_wysiwyg = "true";
defparam \reg_file[6][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N5
dffeas \reg_file[5][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][17] .is_wysiwyg = "true";
defparam \reg_file[5][17] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N3
dffeas \reg_file[4][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][17] .is_wysiwyg = "true";
defparam \reg_file[4][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N4
cycloneive_lcell_comb \Mux46~10 (
// Equation(s):
// \Mux46~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][17]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][17]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][17]~q ),
	.datad(\reg_file[4][17]~q ),
	.cin(gnd),
	.combout(\Mux46~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~10 .lut_mask = 16'hB9A8;
defparam \Mux46~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N0
cycloneive_lcell_comb \Mux46~11 (
// Equation(s):
// \Mux46~11_combout  = (\prif.imemload_id [17] & ((\Mux46~10_combout  & (\reg_file[7][17]~q )) # (!\Mux46~10_combout  & ((\reg_file[6][17]~q ))))) # (!\prif.imemload_id [17] & (((\Mux46~10_combout ))))

	.dataa(\reg_file[7][17]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[6][17]~q ),
	.datad(\Mux46~10_combout ),
	.cin(gnd),
	.combout(\Mux46~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux46~11 .lut_mask = 16'hBBC0;
defparam \Mux46~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N12
cycloneive_lcell_comb \reg_file_nxt[31][21]~88 (
// Equation(s):
// \reg_file_nxt[31][21]~88_combout  = (\Mux143~1_combout  & (((\prif.regwrite_wb [2]) # (\prif.regwrite_wb [0])) # (!Equal8)))

	.dataa(Equal8),
	.datab(prifregwrite_wb_2),
	.datac(Mux143),
	.datad(prifregwrite_wb_0),
	.cin(gnd),
	.combout(\reg_file_nxt[31][21]~88_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][21]~88 .lut_mask = 16'hF0D0;
defparam \reg_file_nxt[31][21]~88 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N24
cycloneive_lcell_comb \reg_file[31][21]~feeder (
// Equation(s):
// \reg_file[31][21]~feeder_combout  = \reg_file_nxt[31][21]~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][21]~88_combout ),
	.cin(gnd),
	.combout(\reg_file[31][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][21]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[31][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N25
dffeas \reg_file[31][21] (
	.clk(!CLK),
	.d(\reg_file[31][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][21] .is_wysiwyg = "true";
defparam \reg_file[31][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N7
dffeas \reg_file[23][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][21] .is_wysiwyg = "true";
defparam \reg_file[23][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N9
dffeas \reg_file[27][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][21] .is_wysiwyg = "true";
defparam \reg_file[27][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N8
cycloneive_lcell_comb \Mux42~7 (
// Equation(s):
// \Mux42~7_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[27][21]~q ))) # (!\prif.imemload_id [19] & (\reg_file[19][21]~q ))))

	.dataa(\reg_file[19][21]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[27][21]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux42~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~7 .lut_mask = 16'hFC22;
defparam \Mux42~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N6
cycloneive_lcell_comb \Mux42~8 (
// Equation(s):
// \Mux42~8_combout  = (\prif.imemload_id [18] & ((\Mux42~7_combout  & (\reg_file[31][21]~q )) # (!\Mux42~7_combout  & ((\reg_file[23][21]~q ))))) # (!\prif.imemload_id [18] & (((\Mux42~7_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[31][21]~q ),
	.datac(\reg_file[23][21]~q ),
	.datad(\Mux42~7_combout ),
	.cin(gnd),
	.combout(\Mux42~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~8 .lut_mask = 16'hDDA0;
defparam \Mux42~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N19
dffeas \reg_file[21][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][21] .is_wysiwyg = "true";
defparam \reg_file[21][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y30_N13
dffeas \reg_file[29][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][21] .is_wysiwyg = "true";
defparam \reg_file[29][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y32_N25
dffeas \reg_file[17][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][21] .is_wysiwyg = "true";
defparam \reg_file[17][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N12
cycloneive_lcell_comb \reg_file[25][21]~feeder (
// Equation(s):
// \reg_file[25][21]~feeder_combout  = \reg_file_nxt[31][21]~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][21]~88_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[25][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][21]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[25][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N13
dffeas \reg_file[25][21] (
	.clk(!CLK),
	.d(\reg_file[25][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][21] .is_wysiwyg = "true";
defparam \reg_file[25][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N24
cycloneive_lcell_comb \Mux42~0 (
// Equation(s):
// \Mux42~0_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[25][21]~q ))) # (!\prif.imemload_id [19] & (\reg_file[17][21]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][21]~q ),
	.datad(\reg_file[25][21]~q ),
	.cin(gnd),
	.combout(\Mux42~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~0 .lut_mask = 16'hDC98;
defparam \Mux42~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N12
cycloneive_lcell_comb \Mux42~1 (
// Equation(s):
// \Mux42~1_combout  = (\prif.imemload_id [18] & ((\Mux42~0_combout  & ((\reg_file[29][21]~q ))) # (!\Mux42~0_combout  & (\reg_file[21][21]~q )))) # (!\prif.imemload_id [18] & (((\Mux42~0_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[21][21]~q ),
	.datac(\reg_file[29][21]~q ),
	.datad(\Mux42~0_combout ),
	.cin(gnd),
	.combout(\Mux42~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~1 .lut_mask = 16'hF588;
defparam \Mux42~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N18
cycloneive_lcell_comb \reg_file[30][21]~feeder (
// Equation(s):
// \reg_file[30][21]~feeder_combout  = \reg_file_nxt[31][21]~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][21]~88_combout ),
	.cin(gnd),
	.combout(\reg_file[30][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[30][21]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[30][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N19
dffeas \reg_file[30][21] (
	.clk(!CLK),
	.d(\reg_file[30][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][21] .is_wysiwyg = "true";
defparam \reg_file[30][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N3
dffeas \reg_file[26][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][21] .is_wysiwyg = "true";
defparam \reg_file[26][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N5
dffeas \reg_file[22][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][21] .is_wysiwyg = "true";
defparam \reg_file[22][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y31_N11
dffeas \reg_file[18][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][21] .is_wysiwyg = "true";
defparam \reg_file[18][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N4
cycloneive_lcell_comb \Mux42~2 (
// Equation(s):
// \Mux42~2_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[22][21]~q )) # (!\prif.imemload_id [18] & ((\reg_file[18][21]~q )))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[22][21]~q ),
	.datad(\reg_file[18][21]~q ),
	.cin(gnd),
	.combout(\Mux42~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~2 .lut_mask = 16'hD9C8;
defparam \Mux42~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N2
cycloneive_lcell_comb \Mux42~3 (
// Equation(s):
// \Mux42~3_combout  = (\prif.imemload_id [19] & ((\Mux42~2_combout  & (\reg_file[30][21]~q )) # (!\Mux42~2_combout  & ((\reg_file[26][21]~q ))))) # (!\prif.imemload_id [19] & (((\Mux42~2_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[30][21]~q ),
	.datac(\reg_file[26][21]~q ),
	.datad(\Mux42~2_combout ),
	.cin(gnd),
	.combout(\Mux42~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~3 .lut_mask = 16'hDDA0;
defparam \Mux42~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N31
dffeas \reg_file[28][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][21] .is_wysiwyg = "true";
defparam \reg_file[28][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N18
cycloneive_lcell_comb \reg_file[20][21]~feeder (
// Equation(s):
// \reg_file[20][21]~feeder_combout  = \reg_file_nxt[31][21]~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][21]~88_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[20][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[20][21]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[20][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N19
dffeas \reg_file[20][21] (
	.clk(!CLK),
	.d(\reg_file[20][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][21] .is_wysiwyg = "true";
defparam \reg_file[20][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N9
dffeas \reg_file[16][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][21] .is_wysiwyg = "true";
defparam \reg_file[16][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N8
cycloneive_lcell_comb \Mux42~4 (
// Equation(s):
// \Mux42~4_combout  = (\prif.imemload_id [18] & ((\reg_file[20][21]~q ) # ((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (((\reg_file[16][21]~q  & !\prif.imemload_id [19]))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[20][21]~q ),
	.datac(\reg_file[16][21]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux42~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~4 .lut_mask = 16'hAAD8;
defparam \Mux42~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N2
cycloneive_lcell_comb \Mux42~5 (
// Equation(s):
// \Mux42~5_combout  = (\prif.imemload_id [19] & ((\Mux42~4_combout  & ((\reg_file[28][21]~q ))) # (!\Mux42~4_combout  & (\reg_file[24][21]~q )))) # (!\prif.imemload_id [19] & (((\Mux42~4_combout ))))

	.dataa(\reg_file[24][21]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[28][21]~q ),
	.datad(\Mux42~4_combout ),
	.cin(gnd),
	.combout(\Mux42~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~5 .lut_mask = 16'hF388;
defparam \Mux42~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N4
cycloneive_lcell_comb \Mux42~6 (
// Equation(s):
// \Mux42~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux42~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & ((\Mux42~5_combout ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux42~3_combout ),
	.datad(\Mux42~5_combout ),
	.cin(gnd),
	.combout(\Mux42~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~6 .lut_mask = 16'hB9A8;
defparam \Mux42~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N13
dffeas \reg_file[15][21] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][21]~88_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][21] .is_wysiwyg = "true";
defparam \reg_file[15][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y31_N25
dffeas \reg_file[14][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][21] .is_wysiwyg = "true";
defparam \reg_file[14][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N25
dffeas \reg_file[13][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][21] .is_wysiwyg = "true";
defparam \reg_file[13][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N7
dffeas \reg_file[12][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][21] .is_wysiwyg = "true";
defparam \reg_file[12][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N24
cycloneive_lcell_comb \Mux42~17 (
// Equation(s):
// \Mux42~17_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[13][21]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[12][21]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[13][21]~q ),
	.datad(\reg_file[12][21]~q ),
	.cin(gnd),
	.combout(\Mux42~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~17 .lut_mask = 16'hB9A8;
defparam \Mux42~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N24
cycloneive_lcell_comb \Mux42~18 (
// Equation(s):
// \Mux42~18_combout  = (\prif.imemload_id [17] & ((\Mux42~17_combout  & (\reg_file[15][21]~q )) # (!\Mux42~17_combout  & ((\reg_file[14][21]~q ))))) # (!\prif.imemload_id [17] & (((\Mux42~17_combout ))))

	.dataa(\reg_file[15][21]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[14][21]~q ),
	.datad(\Mux42~17_combout ),
	.cin(gnd),
	.combout(\Mux42~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~18 .lut_mask = 16'hBBC0;
defparam \Mux42~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N19
dffeas \reg_file[4][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][21] .is_wysiwyg = "true";
defparam \reg_file[4][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N25
dffeas \reg_file[5][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][21] .is_wysiwyg = "true";
defparam \reg_file[5][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N18
cycloneive_lcell_comb \Mux42~10 (
// Equation(s):
// \Mux42~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][21]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & (\reg_file[4][21]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[4][21]~q ),
	.datad(\reg_file[5][21]~q ),
	.cin(gnd),
	.combout(\Mux42~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~10 .lut_mask = 16'hBA98;
defparam \Mux42~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N22
cycloneive_lcell_comb \reg_file[6][21]~feeder (
// Equation(s):
// \reg_file[6][21]~feeder_combout  = \reg_file_nxt[31][21]~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][21]~88_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][21]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N23
dffeas \reg_file[6][21] (
	.clk(!CLK),
	.d(\reg_file[6][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][21] .is_wysiwyg = "true";
defparam \reg_file[6][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y34_N31
dffeas \reg_file[7][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][21] .is_wysiwyg = "true";
defparam \reg_file[7][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N20
cycloneive_lcell_comb \Mux42~11 (
// Equation(s):
// \Mux42~11_combout  = (\prif.imemload_id [17] & ((\Mux42~10_combout  & ((\reg_file[7][21]~q ))) # (!\Mux42~10_combout  & (\reg_file[6][21]~q )))) # (!\prif.imemload_id [17] & (\Mux42~10_combout ))

	.dataa(prifimemload_id_17),
	.datab(\Mux42~10_combout ),
	.datac(\reg_file[6][21]~q ),
	.datad(\reg_file[7][21]~q ),
	.cin(gnd),
	.combout(\Mux42~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~11 .lut_mask = 16'hEC64;
defparam \Mux42~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N27
dffeas \reg_file[1][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][21] .is_wysiwyg = "true";
defparam \reg_file[1][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N0
cycloneive_lcell_comb \reg_file[3][21]~feeder (
// Equation(s):
// \reg_file[3][21]~feeder_combout  = \reg_file_nxt[31][21]~88_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][21]~88_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[3][21]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[3][21]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[3][21]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y33_N1
dffeas \reg_file[3][21] (
	.clk(!CLK),
	.d(\reg_file[3][21]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][21] .is_wysiwyg = "true";
defparam \reg_file[3][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N26
cycloneive_lcell_comb \Mux42~14 (
// Equation(s):
// \Mux42~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][21]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][21]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][21]~q ),
	.datad(\reg_file[3][21]~q ),
	.cin(gnd),
	.combout(\Mux42~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~14 .lut_mask = 16'hC840;
defparam \Mux42~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y34_N1
dffeas \reg_file[2][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][21] .is_wysiwyg = "true";
defparam \reg_file[2][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N8
cycloneive_lcell_comb \Mux42~15 (
// Equation(s):
// \Mux42~15_combout  = (\Mux42~14_combout ) # ((\prif.imemload_id [17] & (!\prif.imemload_id [16] & \reg_file[2][21]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux42~14_combout ),
	.datad(\reg_file[2][21]~q ),
	.cin(gnd),
	.combout(\Mux42~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~15 .lut_mask = 16'hF2F0;
defparam \Mux42~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N25
dffeas \reg_file[11][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][21] .is_wysiwyg = "true";
defparam \reg_file[11][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N3
dffeas \reg_file[8][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][21] .is_wysiwyg = "true";
defparam \reg_file[8][21] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N13
dffeas \reg_file[10][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][21] .is_wysiwyg = "true";
defparam \reg_file[10][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N2
cycloneive_lcell_comb \Mux42~12 (
// Equation(s):
// \Mux42~12_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][21]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][21]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[8][21]~q ),
	.datad(\reg_file[10][21]~q ),
	.cin(gnd),
	.combout(\Mux42~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~12 .lut_mask = 16'hDC98;
defparam \Mux42~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N24
cycloneive_lcell_comb \Mux42~13 (
// Equation(s):
// \Mux42~13_combout  = (\prif.imemload_id [16] & ((\Mux42~12_combout  & ((\reg_file[11][21]~q ))) # (!\Mux42~12_combout  & (\reg_file[9][21]~q )))) # (!\prif.imemload_id [16] & (((\Mux42~12_combout ))))

	.dataa(\reg_file[9][21]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[11][21]~q ),
	.datad(\Mux42~12_combout ),
	.cin(gnd),
	.combout(\Mux42~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~13 .lut_mask = 16'hF388;
defparam \Mux42~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N10
cycloneive_lcell_comb \Mux42~16 (
// Equation(s):
// \Mux42~16_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\Mux42~13_combout ))) # (!\prif.imemload_id [19] & (\Mux42~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux42~15_combout ),
	.datad(\Mux42~13_combout ),
	.cin(gnd),
	.combout(\Mux42~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux42~16 .lut_mask = 16'hDC98;
defparam \Mux42~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N16
cycloneive_lcell_comb \reg_file_nxt[31][20]~89 (
// Equation(s):
// \reg_file_nxt[31][20]~89_combout  = (\Mux144~1_combout  & (((\prif.regwrite_wb [2]) # (\prif.regwrite_wb [0])) # (!Equal8)))

	.dataa(Equal8),
	.datab(prifregwrite_wb_2),
	.datac(Mux144),
	.datad(prifregwrite_wb_0),
	.cin(gnd),
	.combout(\reg_file_nxt[31][20]~89_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][20]~89 .lut_mask = 16'hF0D0;
defparam \reg_file_nxt[31][20]~89 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N28
cycloneive_lcell_comb \reg_file[27][20]~feeder (
// Equation(s):
// \reg_file[27][20]~feeder_combout  = \reg_file_nxt[31][20]~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][20]~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[27][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[27][20]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[27][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N29
dffeas \reg_file[27][20] (
	.clk(!CLK),
	.d(\reg_file[27][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][20] .is_wysiwyg = "true";
defparam \reg_file[27][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N9
dffeas \reg_file[31][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][20] .is_wysiwyg = "true";
defparam \reg_file[31][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N3
dffeas \reg_file[23][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][20] .is_wysiwyg = "true";
defparam \reg_file[23][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N11
dffeas \reg_file[19][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][20] .is_wysiwyg = "true";
defparam \reg_file[19][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N2
cycloneive_lcell_comb \Mux43~7 (
// Equation(s):
// \Mux43~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][20]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][20]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][20]~q ),
	.datad(\reg_file[19][20]~q ),
	.cin(gnd),
	.combout(\Mux43~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~7 .lut_mask = 16'hB9A8;
defparam \Mux43~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N8
cycloneive_lcell_comb \Mux43~8 (
// Equation(s):
// \Mux43~8_combout  = (\prif.imemload_id [19] & ((\Mux43~7_combout  & ((\reg_file[31][20]~q ))) # (!\Mux43~7_combout  & (\reg_file[27][20]~q )))) # (!\prif.imemload_id [19] & (((\Mux43~7_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[27][20]~q ),
	.datac(\reg_file[31][20]~q ),
	.datad(\Mux43~7_combout ),
	.cin(gnd),
	.combout(\Mux43~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~8 .lut_mask = 16'hF588;
defparam \Mux43~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N22
cycloneive_lcell_comb \reg_file[29][20]~feeder (
// Equation(s):
// \reg_file[29][20]~feeder_combout  = \reg_file_nxt[31][20]~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][20]~89_combout ),
	.cin(gnd),
	.combout(\reg_file[29][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][20]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N23
dffeas \reg_file[29][20] (
	.clk(!CLK),
	.d(\reg_file[29][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][20] .is_wysiwyg = "true";
defparam \reg_file[29][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y26_N17
dffeas \reg_file[21][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][20] .is_wysiwyg = "true";
defparam \reg_file[21][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y26_N9
dffeas \reg_file[17][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][20] .is_wysiwyg = "true";
defparam \reg_file[17][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N16
cycloneive_lcell_comb \Mux43~0 (
// Equation(s):
// \Mux43~0_combout  = (\prif.imemload_id [19] & (\prif.imemload_id [18])) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[21][20]~q )) # (!\prif.imemload_id [18] & ((\reg_file[17][20]~q )))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[21][20]~q ),
	.datad(\reg_file[17][20]~q ),
	.cin(gnd),
	.combout(\Mux43~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~0 .lut_mask = 16'hD9C8;
defparam \Mux43~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y26_N23
dffeas \reg_file[25][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][20] .is_wysiwyg = "true";
defparam \reg_file[25][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N22
cycloneive_lcell_comb \Mux43~1 (
// Equation(s):
// \Mux43~1_combout  = (\Mux43~0_combout  & ((\reg_file[29][20]~q ) # ((!\prif.imemload_id [19])))) # (!\Mux43~0_combout  & (((\reg_file[25][20]~q  & \prif.imemload_id [19]))))

	.dataa(\reg_file[29][20]~q ),
	.datab(\Mux43~0_combout ),
	.datac(\reg_file[25][20]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux43~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~1 .lut_mask = 16'hB8CC;
defparam \Mux43~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N29
dffeas \reg_file[20][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][20] .is_wysiwyg = "true";
defparam \reg_file[20][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y33_N15
dffeas \reg_file[28][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][20] .is_wysiwyg = "true";
defparam \reg_file[28][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N24
cycloneive_lcell_comb \reg_file[24][20]~feeder (
// Equation(s):
// \reg_file[24][20]~feeder_combout  = \reg_file_nxt[31][20]~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][20]~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[24][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][20]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[24][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N25
dffeas \reg_file[24][20] (
	.clk(!CLK),
	.d(\reg_file[24][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][20] .is_wysiwyg = "true";
defparam \reg_file[24][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N3
dffeas \reg_file[16][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][20] .is_wysiwyg = "true";
defparam \reg_file[16][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N2
cycloneive_lcell_comb \Mux43~4 (
// Equation(s):
// \Mux43~4_combout  = (\prif.imemload_id [19] & ((\reg_file[24][20]~q ) # ((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (((\reg_file[16][20]~q  & !\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[24][20]~q ),
	.datac(\reg_file[16][20]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux43~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~4 .lut_mask = 16'hAAD8;
defparam \Mux43~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N4
cycloneive_lcell_comb \Mux43~5 (
// Equation(s):
// \Mux43~5_combout  = (\prif.imemload_id [18] & ((\Mux43~4_combout  & ((\reg_file[28][20]~q ))) # (!\Mux43~4_combout  & (\reg_file[20][20]~q )))) # (!\prif.imemload_id [18] & (((\Mux43~4_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[20][20]~q ),
	.datac(\reg_file[28][20]~q ),
	.datad(\Mux43~4_combout ),
	.cin(gnd),
	.combout(\Mux43~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~5 .lut_mask = 16'hF588;
defparam \Mux43~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N21
dffeas \reg_file[22][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][20] .is_wysiwyg = "true";
defparam \reg_file[22][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N11
dffeas \reg_file[30][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][20] .is_wysiwyg = "true";
defparam \reg_file[30][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N20
cycloneive_lcell_comb \Mux43~3 (
// Equation(s):
// \Mux43~3_combout  = (\Mux43~2_combout  & (((\reg_file[30][20]~q )) # (!\prif.imemload_id [18]))) # (!\Mux43~2_combout  & (\prif.imemload_id [18] & (\reg_file[22][20]~q )))

	.dataa(\Mux43~2_combout ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[22][20]~q ),
	.datad(\reg_file[30][20]~q ),
	.cin(gnd),
	.combout(\Mux43~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~3 .lut_mask = 16'hEA62;
defparam \Mux43~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N30
cycloneive_lcell_comb \Mux43~6 (
// Equation(s):
// \Mux43~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux43~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & (\Mux43~5_combout )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux43~5_combout ),
	.datad(\Mux43~3_combout ),
	.cin(gnd),
	.combout(\Mux43~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~6 .lut_mask = 16'hBA98;
defparam \Mux43~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N31
dffeas \reg_file[11][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][20] .is_wysiwyg = "true";
defparam \reg_file[11][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N0
cycloneive_lcell_comb \reg_file[9][20]~feeder (
// Equation(s):
// \reg_file[9][20]~feeder_combout  = \reg_file_nxt[31][20]~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][20]~89_combout ),
	.cin(gnd),
	.combout(\reg_file[9][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[9][20]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[9][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N1
dffeas \reg_file[9][20] (
	.clk(!CLK),
	.d(\reg_file[9][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][20] .is_wysiwyg = "true";
defparam \reg_file[9][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N9
dffeas \reg_file[10][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][20] .is_wysiwyg = "true";
defparam \reg_file[10][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N8
cycloneive_lcell_comb \Mux43~10 (
// Equation(s):
// \Mux43~10_combout  = (\prif.imemload_id [17] & (((\reg_file[10][20]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][20]~q  & ((!\prif.imemload_id [16]))))

	.dataa(\reg_file[8][20]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[10][20]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux43~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~10 .lut_mask = 16'hCCE2;
defparam \Mux43~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N6
cycloneive_lcell_comb \Mux43~11 (
// Equation(s):
// \Mux43~11_combout  = (\prif.imemload_id [16] & ((\Mux43~10_combout  & (\reg_file[11][20]~q )) # (!\Mux43~10_combout  & ((\reg_file[9][20]~q ))))) # (!\prif.imemload_id [16] & (((\Mux43~10_combout ))))

	.dataa(\reg_file[11][20]~q ),
	.datab(\reg_file[9][20]~q ),
	.datac(prifimemload_id_16),
	.datad(\Mux43~10_combout ),
	.cin(gnd),
	.combout(\Mux43~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~11 .lut_mask = 16'hAFC0;
defparam \Mux43~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N17
dffeas \reg_file[15][20] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][20]~89_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][20] .is_wysiwyg = "true";
defparam \reg_file[15][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y31_N11
dffeas \reg_file[14][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][20] .is_wysiwyg = "true";
defparam \reg_file[14][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y31_N21
dffeas \reg_file[13][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][20] .is_wysiwyg = "true";
defparam \reg_file[13][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N20
cycloneive_lcell_comb \Mux43~17 (
// Equation(s):
// \Mux43~17_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][20]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][20]~q ))))

	.dataa(\reg_file[12][20]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[13][20]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux43~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~17 .lut_mask = 16'hFC22;
defparam \Mux43~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N10
cycloneive_lcell_comb \Mux43~18 (
// Equation(s):
// \Mux43~18_combout  = (\prif.imemload_id [17] & ((\Mux43~17_combout  & (\reg_file[15][20]~q )) # (!\Mux43~17_combout  & ((\reg_file[14][20]~q ))))) # (!\prif.imemload_id [17] & (((\Mux43~17_combout ))))

	.dataa(\reg_file[15][20]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[14][20]~q ),
	.datad(\Mux43~17_combout ),
	.cin(gnd),
	.combout(\Mux43~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~18 .lut_mask = 16'hBBC0;
defparam \Mux43~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N13
dffeas \reg_file[5][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][20] .is_wysiwyg = "true";
defparam \reg_file[5][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N7
dffeas \reg_file[4][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][20] .is_wysiwyg = "true";
defparam \reg_file[4][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N12
cycloneive_lcell_comb \Mux43~12 (
// Equation(s):
// \Mux43~12_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][20]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][20]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][20]~q ),
	.datad(\reg_file[4][20]~q ),
	.cin(gnd),
	.combout(\Mux43~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~12 .lut_mask = 16'hB9A8;
defparam \Mux43~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N5
dffeas \reg_file[7][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][20] .is_wysiwyg = "true";
defparam \reg_file[7][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N4
cycloneive_lcell_comb \Mux43~13 (
// Equation(s):
// \Mux43~13_combout  = (\Mux43~12_combout  & (((\reg_file[7][20]~q ) # (!\prif.imemload_id [17])))) # (!\Mux43~12_combout  & (\reg_file[6][20]~q  & ((\prif.imemload_id [17]))))

	.dataa(\reg_file[6][20]~q ),
	.datab(\Mux43~12_combout ),
	.datac(\reg_file[7][20]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux43~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~13 .lut_mask = 16'hE2CC;
defparam \Mux43~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N17
dffeas \reg_file[2][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][20] .is_wysiwyg = "true";
defparam \reg_file[2][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N5
dffeas \reg_file[3][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][20] .is_wysiwyg = "true";
defparam \reg_file[3][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N2
cycloneive_lcell_comb \reg_file[1][20]~feeder (
// Equation(s):
// \reg_file[1][20]~feeder_combout  = \reg_file_nxt[31][20]~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][20]~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[1][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[1][20]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[1][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y33_N3
dffeas \reg_file[1][20] (
	.clk(!CLK),
	.d(\reg_file[1][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][20] .is_wysiwyg = "true";
defparam \reg_file[1][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N4
cycloneive_lcell_comb \Mux43~14 (
// Equation(s):
// \Mux43~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][20]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][20]~q )))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[3][20]~q ),
	.datad(\reg_file[1][20]~q ),
	.cin(gnd),
	.combout(\Mux43~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~14 .lut_mask = 16'hC480;
defparam \Mux43~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N12
cycloneive_lcell_comb \Mux43~15 (
// Equation(s):
// \Mux43~15_combout  = (\Mux43~14_combout ) # ((!\prif.imemload_id [16] & (\reg_file[2][20]~q  & \prif.imemload_id [17])))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[2][20]~q ),
	.datac(\Mux43~14_combout ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux43~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~15 .lut_mask = 16'hF4F0;
defparam \Mux43~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N18
cycloneive_lcell_comb \Mux43~16 (
// Equation(s):
// \Mux43~16_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\Mux43~13_combout )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\Mux43~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux43~13_combout ),
	.datad(\Mux43~15_combout ),
	.cin(gnd),
	.combout(\Mux43~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux43~16 .lut_mask = 16'hB9A8;
defparam \Mux43~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N20
cycloneive_lcell_comb \reg_file_nxt[31][28]~90 (
// Equation(s):
// \reg_file_nxt[31][28]~90_combout  = (\Mux136~1_combout  & (((\prif.regwrite_wb [2]) # (\prif.regwrite_wb [0])) # (!Equal8)))

	.dataa(Equal8),
	.datab(prifregwrite_wb_2),
	.datac(Mux136),
	.datad(prifregwrite_wb_0),
	.cin(gnd),
	.combout(\reg_file_nxt[31][28]~90_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][28]~90 .lut_mask = 16'hF0D0;
defparam \reg_file_nxt[31][28]~90 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N4
cycloneive_lcell_comb \reg_file[29][28]~feeder (
// Equation(s):
// \reg_file[29][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][28]~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][28]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N5
dffeas \reg_file[29][28] (
	.clk(!CLK),
	.d(\reg_file[29][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][28] .is_wysiwyg = "true";
defparam \reg_file[29][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N4
cycloneive_lcell_comb \reg_file[17][28]~feeder (
// Equation(s):
// \reg_file[17][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][28]~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[17][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[17][28]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[17][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N5
dffeas \reg_file[17][28] (
	.clk(!CLK),
	.d(\reg_file[17][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][28] .is_wysiwyg = "true";
defparam \reg_file[17][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N31
dffeas \reg_file[21][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][28] .is_wysiwyg = "true";
defparam \reg_file[21][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N30
cycloneive_lcell_comb \Mux35~0 (
// Equation(s):
// \Mux35~0_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[21][28]~q ))) # (!\prif.imemload_id [18] & (\reg_file[17][28]~q ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[17][28]~q ),
	.datac(\reg_file[21][28]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux35~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~0 .lut_mask = 16'hFA44;
defparam \Mux35~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N28
cycloneive_lcell_comb \reg_file[25][28]~feeder (
// Equation(s):
// \reg_file[25][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][28]~90_combout ),
	.cin(gnd),
	.combout(\reg_file[25][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][28]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[25][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N29
dffeas \reg_file[25][28] (
	.clk(!CLK),
	.d(\reg_file[25][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][28] .is_wysiwyg = "true";
defparam \reg_file[25][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N18
cycloneive_lcell_comb \Mux35~1 (
// Equation(s):
// \Mux35~1_combout  = (\prif.imemload_id [19] & ((\Mux35~0_combout  & (\reg_file[29][28]~q )) # (!\Mux35~0_combout  & ((\reg_file[25][28]~q ))))) # (!\prif.imemload_id [19] & (((\Mux35~0_combout ))))

	.dataa(\reg_file[29][28]~q ),
	.datab(prifimemload_id_19),
	.datac(\Mux35~0_combout ),
	.datad(\reg_file[25][28]~q ),
	.cin(gnd),
	.combout(\Mux35~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~1 .lut_mask = 16'hBCB0;
defparam \Mux35~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N15
dffeas \reg_file[30][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][28] .is_wysiwyg = "true";
defparam \reg_file[30][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N20
cycloneive_lcell_comb \reg_file[22][28]~feeder (
// Equation(s):
// \reg_file[22][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][28]~90_combout ),
	.cin(gnd),
	.combout(\reg_file[22][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][28]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[22][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N21
dffeas \reg_file[22][28] (
	.clk(!CLK),
	.d(\reg_file[22][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][28] .is_wysiwyg = "true";
defparam \reg_file[22][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N6
cycloneive_lcell_comb \Mux35~3 (
// Equation(s):
// \Mux35~3_combout  = (\Mux35~2_combout  & ((\reg_file[30][28]~q ) # ((!\prif.imemload_id [18])))) # (!\Mux35~2_combout  & (((\prif.imemload_id [18] & \reg_file[22][28]~q ))))

	.dataa(\Mux35~2_combout ),
	.datab(\reg_file[30][28]~q ),
	.datac(prifimemload_id_18),
	.datad(\reg_file[22][28]~q ),
	.cin(gnd),
	.combout(\Mux35~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~3 .lut_mask = 16'hDA8A;
defparam \Mux35~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N19
dffeas \reg_file[28][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][28] .is_wysiwyg = "true";
defparam \reg_file[28][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N11
dffeas \reg_file[20][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][28] .is_wysiwyg = "true";
defparam \reg_file[20][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N28
cycloneive_lcell_comb \reg_file[24][28]~feeder (
// Equation(s):
// \reg_file[24][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][28]~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[24][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][28]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[24][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N29
dffeas \reg_file[24][28] (
	.clk(!CLK),
	.d(\reg_file[24][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][28] .is_wysiwyg = "true";
defparam \reg_file[24][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N21
dffeas \reg_file[16][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][28] .is_wysiwyg = "true";
defparam \reg_file[16][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N20
cycloneive_lcell_comb \Mux35~4 (
// Equation(s):
// \Mux35~4_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[24][28]~q )) # (!\prif.imemload_id [19] & ((\reg_file[16][28]~q )))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[24][28]~q ),
	.datac(\reg_file[16][28]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux35~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~4 .lut_mask = 16'hEE50;
defparam \Mux35~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N28
cycloneive_lcell_comb \Mux35~5 (
// Equation(s):
// \Mux35~5_combout  = (\prif.imemload_id [18] & ((\Mux35~4_combout  & (\reg_file[28][28]~q )) # (!\Mux35~4_combout  & ((\reg_file[20][28]~q ))))) # (!\prif.imemload_id [18] & (((\Mux35~4_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[28][28]~q ),
	.datac(\reg_file[20][28]~q ),
	.datad(\Mux35~4_combout ),
	.cin(gnd),
	.combout(\Mux35~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~5 .lut_mask = 16'hDDA0;
defparam \Mux35~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N22
cycloneive_lcell_comb \Mux35~6 (
// Equation(s):
// \Mux35~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux35~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & ((\Mux35~5_combout ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux35~3_combout ),
	.datad(\Mux35~5_combout ),
	.cin(gnd),
	.combout(\Mux35~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~6 .lut_mask = 16'hB9A8;
defparam \Mux35~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y29_N31
dffeas \reg_file[23][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][28] .is_wysiwyg = "true";
defparam \reg_file[23][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N15
dffeas \reg_file[19][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][28] .is_wysiwyg = "true";
defparam \reg_file[19][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N30
cycloneive_lcell_comb \Mux35~7 (
// Equation(s):
// \Mux35~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][28]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][28]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][28]~q ),
	.datad(\reg_file[19][28]~q ),
	.cin(gnd),
	.combout(\Mux35~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~7 .lut_mask = 16'hB9A8;
defparam \Mux35~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N29
dffeas \reg_file[27][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][28] .is_wysiwyg = "true";
defparam \reg_file[27][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N1
dffeas \reg_file[31][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][28] .is_wysiwyg = "true";
defparam \reg_file[31][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N28
cycloneive_lcell_comb \Mux35~8 (
// Equation(s):
// \Mux35~8_combout  = (\prif.imemload_id [19] & ((\Mux35~7_combout  & ((\reg_file[31][28]~q ))) # (!\Mux35~7_combout  & (\reg_file[27][28]~q )))) # (!\prif.imemload_id [19] & (\Mux35~7_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux35~7_combout ),
	.datac(\reg_file[27][28]~q ),
	.datad(\reg_file[31][28]~q ),
	.cin(gnd),
	.combout(\Mux35~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~8 .lut_mask = 16'hEC64;
defparam \Mux35~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N18
cycloneive_lcell_comb \reg_file[9][28]~feeder (
// Equation(s):
// \reg_file[9][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][28]~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[9][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[9][28]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[9][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N19
dffeas \reg_file[9][28] (
	.clk(!CLK),
	.d(\reg_file[9][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][28] .is_wysiwyg = "true";
defparam \reg_file[9][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N12
cycloneive_lcell_comb \reg_file[11][28]~feeder (
// Equation(s):
// \reg_file[11][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][28]~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[11][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[11][28]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[11][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N13
dffeas \reg_file[11][28] (
	.clk(!CLK),
	.d(\reg_file[11][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][28] .is_wysiwyg = "true";
defparam \reg_file[11][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N5
dffeas \reg_file[10][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][28] .is_wysiwyg = "true";
defparam \reg_file[10][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N4
cycloneive_lcell_comb \Mux35~10 (
// Equation(s):
// \Mux35~10_combout  = (\prif.imemload_id [17] & (((\reg_file[10][28]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][28]~q  & ((!\prif.imemload_id [16]))))

	.dataa(\reg_file[8][28]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[10][28]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux35~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~10 .lut_mask = 16'hCCE2;
defparam \Mux35~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N12
cycloneive_lcell_comb \Mux35~11 (
// Equation(s):
// \Mux35~11_combout  = (\Mux35~10_combout  & (((\reg_file[11][28]~q ) # (!\prif.imemload_id [16])))) # (!\Mux35~10_combout  & (\reg_file[9][28]~q  & ((\prif.imemload_id [16]))))

	.dataa(\reg_file[9][28]~q ),
	.datab(\reg_file[11][28]~q ),
	.datac(\Mux35~10_combout ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux35~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~11 .lut_mask = 16'hCAF0;
defparam \Mux35~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N12
cycloneive_lcell_comb \reg_file[14][28]~feeder (
// Equation(s):
// \reg_file[14][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][28]~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[14][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][28]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[14][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N13
dffeas \reg_file[14][28] (
	.clk(!CLK),
	.d(\reg_file[14][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][28] .is_wysiwyg = "true";
defparam \reg_file[14][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N17
dffeas \reg_file[13][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][28] .is_wysiwyg = "true";
defparam \reg_file[13][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N16
cycloneive_lcell_comb \Mux35~17 (
// Equation(s):
// \Mux35~17_combout  = (\prif.imemload_id [16] & (((\reg_file[13][28]~q ) # (\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & (\reg_file[12][28]~q  & ((!\prif.imemload_id [17]))))

	.dataa(\reg_file[12][28]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[13][28]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux35~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~17 .lut_mask = 16'hCCE2;
defparam \Mux35~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N21
dffeas \reg_file[15][28] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][28]~90_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][28] .is_wysiwyg = "true";
defparam \reg_file[15][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N6
cycloneive_lcell_comb \Mux35~18 (
// Equation(s):
// \Mux35~18_combout  = (\Mux35~17_combout  & (((\reg_file[15][28]~q ) # (!\prif.imemload_id [17])))) # (!\Mux35~17_combout  & (\reg_file[14][28]~q  & (\prif.imemload_id [17])))

	.dataa(\reg_file[14][28]~q ),
	.datab(\Mux35~17_combout ),
	.datac(prifimemload_id_17),
	.datad(\reg_file[15][28]~q ),
	.cin(gnd),
	.combout(\Mux35~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~18 .lut_mask = 16'hEC2C;
defparam \Mux35~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N18
cycloneive_lcell_comb \reg_file[2][28]~feeder (
// Equation(s):
// \reg_file[2][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][28]~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[2][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][28]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[2][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N19
dffeas \reg_file[2][28] (
	.clk(!CLK),
	.d(\reg_file[2][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][28] .is_wysiwyg = "true";
defparam \reg_file[2][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N14
cycloneive_lcell_comb \reg_file[1][28]~feeder (
// Equation(s):
// \reg_file[1][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][28]~90_combout ),
	.cin(gnd),
	.combout(\reg_file[1][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[1][28]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[1][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y34_N15
dffeas \reg_file[1][28] (
	.clk(!CLK),
	.d(\reg_file[1][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][28] .is_wysiwyg = "true";
defparam \reg_file[1][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y34_N29
dffeas \reg_file[3][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][28] .is_wysiwyg = "true";
defparam \reg_file[3][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N28
cycloneive_lcell_comb \Mux35~14 (
// Equation(s):
// \Mux35~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][28]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][28]~q ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[1][28]~q ),
	.datac(\reg_file[3][28]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux35~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~14 .lut_mask = 16'hA088;
defparam \Mux35~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N24
cycloneive_lcell_comb \Mux35~15 (
// Equation(s):
// \Mux35~15_combout  = (\Mux35~14_combout ) # ((\prif.imemload_id [17] & (!\prif.imemload_id [16] & \reg_file[2][28]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[2][28]~q ),
	.datad(\Mux35~14_combout ),
	.cin(gnd),
	.combout(\Mux35~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~15 .lut_mask = 16'hFF20;
defparam \Mux35~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N12
cycloneive_lcell_comb \reg_file[7][28]~feeder (
// Equation(s):
// \reg_file[7][28]~feeder_combout  = \reg_file_nxt[31][28]~90_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][28]~90_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[7][28]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[7][28]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[7][28]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N13
dffeas \reg_file[7][28] (
	.clk(!CLK),
	.d(\reg_file[7][28]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][28] .is_wysiwyg = "true";
defparam \reg_file[7][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N19
dffeas \reg_file[6][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][28] .is_wysiwyg = "true";
defparam \reg_file[6][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N18
cycloneive_lcell_comb \Mux35~13 (
// Equation(s):
// \Mux35~13_combout  = (\Mux35~12_combout  & (((\reg_file[7][28]~q )) # (!\prif.imemload_id [17]))) # (!\Mux35~12_combout  & (\prif.imemload_id [17] & ((\reg_file[6][28]~q ))))

	.dataa(\Mux35~12_combout ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[7][28]~q ),
	.datad(\reg_file[6][28]~q ),
	.cin(gnd),
	.combout(\Mux35~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~13 .lut_mask = 16'hE6A2;
defparam \Mux35~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y33_N28
cycloneive_lcell_comb \Mux35~16 (
// Equation(s):
// \Mux35~16_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\Mux35~13_combout ))) # (!\prif.imemload_id [18] & (\Mux35~15_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\Mux35~15_combout ),
	.datac(\Mux35~13_combout ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux35~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux35~16 .lut_mask = 16'hFA44;
defparam \Mux35~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N30
cycloneive_lcell_comb \reg_file_nxt[31][26]~91 (
// Equation(s):
// \reg_file_nxt[31][26]~91_combout  = (\Mux138~1_combout  & (((\prif.regwrite_wb [2]) # (\prif.regwrite_wb [0])) # (!Equal8)))

	.dataa(Equal8),
	.datab(prifregwrite_wb_2),
	.datac(Mux138),
	.datad(prifregwrite_wb_0),
	.cin(gnd),
	.combout(\reg_file_nxt[31][26]~91_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][26]~91 .lut_mask = 16'hF0D0;
defparam \reg_file_nxt[31][26]~91 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N26
cycloneive_lcell_comb \reg_file[22][26]~feeder (
// Equation(s):
// \reg_file[22][26]~feeder_combout  = \reg_file_nxt[31][26]~91_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][26]~91_combout ),
	.cin(gnd),
	.combout(\reg_file[22][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][26]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[22][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N27
dffeas \reg_file[22][26] (
	.clk(!CLK),
	.d(\reg_file[22][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][26] .is_wysiwyg = "true";
defparam \reg_file[22][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y31_N5
dffeas \reg_file[30][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][26] .is_wysiwyg = "true";
defparam \reg_file[30][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N4
cycloneive_lcell_comb \Mux37~3 (
// Equation(s):
// \Mux37~3_combout  = (\Mux37~2_combout  & (((\reg_file[30][26]~q ) # (!\prif.imemload_id [18])))) # (!\Mux37~2_combout  & (\reg_file[22][26]~q  & ((\prif.imemload_id [18]))))

	.dataa(\Mux37~2_combout ),
	.datab(\reg_file[22][26]~q ),
	.datac(\reg_file[30][26]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux37~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~3 .lut_mask = 16'hE4AA;
defparam \Mux37~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N1
dffeas \reg_file[20][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][26] .is_wysiwyg = "true";
defparam \reg_file[20][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N15
dffeas \reg_file[28][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][26] .is_wysiwyg = "true";
defparam \reg_file[28][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N14
cycloneive_lcell_comb \Mux37~5 (
// Equation(s):
// \Mux37~5_combout  = (\Mux37~4_combout  & (((\reg_file[28][26]~q ) # (!\prif.imemload_id [18])))) # (!\Mux37~4_combout  & (\reg_file[20][26]~q  & ((\prif.imemload_id [18]))))

	.dataa(\Mux37~4_combout ),
	.datab(\reg_file[20][26]~q ),
	.datac(\reg_file[28][26]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux37~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~5 .lut_mask = 16'hE4AA;
defparam \Mux37~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N12
cycloneive_lcell_comb \Mux37~6 (
// Equation(s):
// \Mux37~6_combout  = (\prif.imemload_id [16] & (((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\Mux37~3_combout )) # (!\prif.imemload_id [17] & ((\Mux37~5_combout )))))

	.dataa(\Mux37~3_combout ),
	.datab(\Mux37~5_combout ),
	.datac(prifimemload_id_16),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux37~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~6 .lut_mask = 16'hFA0C;
defparam \Mux37~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N30
cycloneive_lcell_comb \reg_file[29][26]~feeder (
// Equation(s):
// \reg_file[29][26]~feeder_combout  = \reg_file_nxt[31][26]~91_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][26]~91_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][26]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N31
dffeas \reg_file[29][26] (
	.clk(!CLK),
	.d(\reg_file[29][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][26] .is_wysiwyg = "true";
defparam \reg_file[29][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y30_N1
dffeas \reg_file[25][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][26] .is_wysiwyg = "true";
defparam \reg_file[25][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N3
dffeas \reg_file[17][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][26] .is_wysiwyg = "true";
defparam \reg_file[17][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N9
dffeas \reg_file[21][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][26] .is_wysiwyg = "true";
defparam \reg_file[21][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N8
cycloneive_lcell_comb \Mux37~0 (
// Equation(s):
// \Mux37~0_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[21][26]~q ))) # (!\prif.imemload_id [18] & (\reg_file[17][26]~q ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[17][26]~q ),
	.datac(\reg_file[21][26]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux37~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~0 .lut_mask = 16'hFA44;
defparam \Mux37~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N0
cycloneive_lcell_comb \Mux37~1 (
// Equation(s):
// \Mux37~1_combout  = (\prif.imemload_id [19] & ((\Mux37~0_combout  & (\reg_file[29][26]~q )) # (!\Mux37~0_combout  & ((\reg_file[25][26]~q ))))) # (!\prif.imemload_id [19] & (((\Mux37~0_combout ))))

	.dataa(\reg_file[29][26]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[25][26]~q ),
	.datad(\Mux37~0_combout ),
	.cin(gnd),
	.combout(\Mux37~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~1 .lut_mask = 16'hBBC0;
defparam \Mux37~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y27_N13
dffeas \reg_file[31][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][26] .is_wysiwyg = "true";
defparam \reg_file[31][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y27_N5
dffeas \reg_file[27][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][26] .is_wysiwyg = "true";
defparam \reg_file[27][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N17
dffeas \reg_file[23][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][26] .is_wysiwyg = "true";
defparam \reg_file[23][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N27
dffeas \reg_file[19][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][26] .is_wysiwyg = "true";
defparam \reg_file[19][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N16
cycloneive_lcell_comb \Mux37~7 (
// Equation(s):
// \Mux37~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][26]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][26]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][26]~q ),
	.datad(\reg_file[19][26]~q ),
	.cin(gnd),
	.combout(\Mux37~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~7 .lut_mask = 16'hB9A8;
defparam \Mux37~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N4
cycloneive_lcell_comb \Mux37~8 (
// Equation(s):
// \Mux37~8_combout  = (\prif.imemload_id [19] & ((\Mux37~7_combout  & (\reg_file[31][26]~q )) # (!\Mux37~7_combout  & ((\reg_file[27][26]~q ))))) # (!\prif.imemload_id [19] & (((\Mux37~7_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[31][26]~q ),
	.datac(\reg_file[27][26]~q ),
	.datad(\Mux37~7_combout ),
	.cin(gnd),
	.combout(\Mux37~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~8 .lut_mask = 16'hDDA0;
defparam \Mux37~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N29
dffeas \reg_file[10][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][26] .is_wysiwyg = "true";
defparam \reg_file[10][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N28
cycloneive_lcell_comb \Mux37~10 (
// Equation(s):
// \Mux37~10_combout  = (\prif.imemload_id [17] & (((\reg_file[10][26]~q ) # (\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & (\reg_file[8][26]~q  & ((!\prif.imemload_id [16]))))

	.dataa(\reg_file[8][26]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[10][26]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux37~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~10 .lut_mask = 16'hCCE2;
defparam \Mux37~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y31_N1
dffeas \reg_file[9][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][26] .is_wysiwyg = "true";
defparam \reg_file[9][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N16
cycloneive_lcell_comb \reg_file[11][26]~feeder (
// Equation(s):
// \reg_file[11][26]~feeder_combout  = \reg_file_nxt[31][26]~91_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][26]~91_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[11][26]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[11][26]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[11][26]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N17
dffeas \reg_file[11][26] (
	.clk(!CLK),
	.d(\reg_file[11][26]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][26] .is_wysiwyg = "true";
defparam \reg_file[11][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N0
cycloneive_lcell_comb \Mux37~11 (
// Equation(s):
// \Mux37~11_combout  = (\prif.imemload_id [16] & ((\Mux37~10_combout  & ((\reg_file[11][26]~q ))) # (!\Mux37~10_combout  & (\reg_file[9][26]~q )))) # (!\prif.imemload_id [16] & (\Mux37~10_combout ))

	.dataa(prifimemload_id_16),
	.datab(\Mux37~10_combout ),
	.datac(\reg_file[9][26]~q ),
	.datad(\reg_file[11][26]~q ),
	.cin(gnd),
	.combout(\Mux37~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~11 .lut_mask = 16'hEC64;
defparam \Mux37~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y31_N31
dffeas \reg_file[15][26] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][26]~91_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][26] .is_wysiwyg = "true";
defparam \reg_file[15][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N21
dffeas \reg_file[14][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][26] .is_wysiwyg = "true";
defparam \reg_file[14][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N13
dffeas \reg_file[13][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][26] .is_wysiwyg = "true";
defparam \reg_file[13][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N12
cycloneive_lcell_comb \Mux37~17 (
// Equation(s):
// \Mux37~17_combout  = (\prif.imemload_id [16] & (((\reg_file[13][26]~q ) # (\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & (\reg_file[12][26]~q  & ((!\prif.imemload_id [17]))))

	.dataa(\reg_file[12][26]~q ),
	.datab(prifimemload_id_16),
	.datac(\reg_file[13][26]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux37~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~17 .lut_mask = 16'hCCE2;
defparam \Mux37~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N20
cycloneive_lcell_comb \Mux37~18 (
// Equation(s):
// \Mux37~18_combout  = (\prif.imemload_id [17] & ((\Mux37~17_combout  & (\reg_file[15][26]~q )) # (!\Mux37~17_combout  & ((\reg_file[14][26]~q ))))) # (!\prif.imemload_id [17] & (((\Mux37~17_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[15][26]~q ),
	.datac(\reg_file[14][26]~q ),
	.datad(\Mux37~17_combout ),
	.cin(gnd),
	.combout(\Mux37~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~18 .lut_mask = 16'hDDA0;
defparam \Mux37~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N9
dffeas \reg_file[6][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][26] .is_wysiwyg = "true";
defparam \reg_file[6][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N7
dffeas \reg_file[7][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][26] .is_wysiwyg = "true";
defparam \reg_file[7][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N5
dffeas \reg_file[5][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][26] .is_wysiwyg = "true";
defparam \reg_file[5][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N4
cycloneive_lcell_comb \Mux37~12 (
// Equation(s):
// \Mux37~12_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[5][26]~q ))) # (!\prif.imemload_id [16] & (\reg_file[4][26]~q ))))

	.dataa(\reg_file[4][26]~q ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][26]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux37~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~12 .lut_mask = 16'hFC22;
defparam \Mux37~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N6
cycloneive_lcell_comb \Mux37~13 (
// Equation(s):
// \Mux37~13_combout  = (\prif.imemload_id [17] & ((\Mux37~12_combout  & ((\reg_file[7][26]~q ))) # (!\Mux37~12_combout  & (\reg_file[6][26]~q )))) # (!\prif.imemload_id [17] & (((\Mux37~12_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[6][26]~q ),
	.datac(\reg_file[7][26]~q ),
	.datad(\Mux37~12_combout ),
	.cin(gnd),
	.combout(\Mux37~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~13 .lut_mask = 16'hF588;
defparam \Mux37~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N17
dffeas \reg_file[1][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][26] .is_wysiwyg = "true";
defparam \reg_file[1][26] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N7
dffeas \reg_file[3][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][26] .is_wysiwyg = "true";
defparam \reg_file[3][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N16
cycloneive_lcell_comb \Mux37~14 (
// Equation(s):
// \Mux37~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][26]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][26]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][26]~q ),
	.datad(\reg_file[3][26]~q ),
	.cin(gnd),
	.combout(\Mux37~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~14 .lut_mask = 16'hC840;
defparam \Mux37~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N15
dffeas \reg_file[2][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][26] .is_wysiwyg = "true";
defparam \reg_file[2][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N28
cycloneive_lcell_comb \Mux37~15 (
// Equation(s):
// \Mux37~15_combout  = (\Mux37~14_combout ) # ((\prif.imemload_id [17] & (!\prif.imemload_id [16] & \reg_file[2][26]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux37~14_combout ),
	.datad(\reg_file[2][26]~q ),
	.cin(gnd),
	.combout(\Mux37~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~15 .lut_mask = 16'hF2F0;
defparam \Mux37~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y32_N6
cycloneive_lcell_comb \Mux37~16 (
// Equation(s):
// \Mux37~16_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\Mux37~13_combout )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\Mux37~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux37~13_combout ),
	.datad(\Mux37~15_combout ),
	.cin(gnd),
	.combout(\Mux37~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux37~16 .lut_mask = 16'hB9A8;
defparam \Mux37~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N0
cycloneive_lcell_comb \reg_file_nxt[31][8]~92 (
// Equation(s):
// \reg_file_nxt[31][8]~92_combout  = (\Mux156~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(prifregwrite_wb_0),
	.datac(Mux156),
	.datad(Equal8),
	.cin(gnd),
	.combout(\reg_file_nxt[31][8]~92_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][8]~92 .lut_mask = 16'hE0F0;
defparam \reg_file_nxt[31][8]~92 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N11
dffeas \reg_file[29][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][8] .is_wysiwyg = "true";
defparam \reg_file[29][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N15
dffeas \reg_file[17][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][8] .is_wysiwyg = "true";
defparam \reg_file[17][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N4
cycloneive_lcell_comb \Mux55~0 (
// Equation(s):
// \Mux55~0_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & (\reg_file[21][8]~q )) # (!\prif.imemload_id [18] & ((\reg_file[17][8]~q )))))

	.dataa(\reg_file[21][8]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[17][8]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux55~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~0 .lut_mask = 16'hEE30;
defparam \Mux55~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N10
cycloneive_lcell_comb \reg_file[25][8]~feeder (
// Equation(s):
// \reg_file[25][8]~feeder_combout  = \reg_file_nxt[31][8]~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][8]~92_combout ),
	.cin(gnd),
	.combout(\reg_file[25][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][8]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[25][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N11
dffeas \reg_file[25][8] (
	.clk(!CLK),
	.d(\reg_file[25][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][8] .is_wysiwyg = "true";
defparam \reg_file[25][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N18
cycloneive_lcell_comb \Mux55~1 (
// Equation(s):
// \Mux55~1_combout  = (\prif.imemload_id [19] & ((\Mux55~0_combout  & (\reg_file[29][8]~q )) # (!\Mux55~0_combout  & ((\reg_file[25][8]~q ))))) # (!\prif.imemload_id [19] & (((\Mux55~0_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[29][8]~q ),
	.datac(\Mux55~0_combout ),
	.datad(\reg_file[25][8]~q ),
	.cin(gnd),
	.combout(\Mux55~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~1 .lut_mask = 16'hDAD0;
defparam \Mux55~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y27_N3
dffeas \reg_file[23][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][8] .is_wysiwyg = "true";
defparam \reg_file[23][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N19
dffeas \reg_file[19][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][8] .is_wysiwyg = "true";
defparam \reg_file[19][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y27_N2
cycloneive_lcell_comb \Mux55~7 (
// Equation(s):
// \Mux55~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][8]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][8]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][8]~q ),
	.datad(\reg_file[19][8]~q ),
	.cin(gnd),
	.combout(\Mux55~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~7 .lut_mask = 16'hB9A8;
defparam \Mux55~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y28_N17
dffeas \reg_file[27][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][8] .is_wysiwyg = "true";
defparam \reg_file[27][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N12
cycloneive_lcell_comb \reg_file[31][8]~feeder (
// Equation(s):
// \reg_file[31][8]~feeder_combout  = \reg_file_nxt[31][8]~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][8]~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[31][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[31][8]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[31][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y26_N13
dffeas \reg_file[31][8] (
	.clk(!CLK),
	.d(\reg_file[31][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][8] .is_wysiwyg = "true";
defparam \reg_file[31][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N16
cycloneive_lcell_comb \Mux55~8 (
// Equation(s):
// \Mux55~8_combout  = (\Mux55~7_combout  & (((\reg_file[31][8]~q )) # (!\prif.imemload_id [19]))) # (!\Mux55~7_combout  & (\prif.imemload_id [19] & (\reg_file[27][8]~q )))

	.dataa(\Mux55~7_combout ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][8]~q ),
	.datad(\reg_file[31][8]~q ),
	.cin(gnd),
	.combout(\Mux55~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~8 .lut_mask = 16'hEA62;
defparam \Mux55~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N5
dffeas \reg_file[20][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][8] .is_wysiwyg = "true";
defparam \reg_file[20][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y32_N31
dffeas \reg_file[28][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][8] .is_wysiwyg = "true";
defparam \reg_file[28][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N23
dffeas \reg_file[16][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][8] .is_wysiwyg = "true";
defparam \reg_file[16][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N26
cycloneive_lcell_comb \reg_file[24][8]~feeder (
// Equation(s):
// \reg_file[24][8]~feeder_combout  = \reg_file_nxt[31][8]~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][8]~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[24][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][8]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[24][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N27
dffeas \reg_file[24][8] (
	.clk(!CLK),
	.d(\reg_file[24][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][8] .is_wysiwyg = "true";
defparam \reg_file[24][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N22
cycloneive_lcell_comb \Mux55~4 (
// Equation(s):
// \Mux55~4_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[24][8]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & (\reg_file[16][8]~q )))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[16][8]~q ),
	.datad(\reg_file[24][8]~q ),
	.cin(gnd),
	.combout(\Mux55~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~4 .lut_mask = 16'hBA98;
defparam \Mux55~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N12
cycloneive_lcell_comb \Mux55~5 (
// Equation(s):
// \Mux55~5_combout  = (\prif.imemload_id [18] & ((\Mux55~4_combout  & ((\reg_file[28][8]~q ))) # (!\Mux55~4_combout  & (\reg_file[20][8]~q )))) # (!\prif.imemload_id [18] & (((\Mux55~4_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[20][8]~q ),
	.datac(\reg_file[28][8]~q ),
	.datad(\Mux55~4_combout ),
	.cin(gnd),
	.combout(\Mux55~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~5 .lut_mask = 16'hF588;
defparam \Mux55~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N29
dffeas \reg_file[18][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][8] .is_wysiwyg = "true";
defparam \reg_file[18][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N19
dffeas \reg_file[26][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][8] .is_wysiwyg = "true";
defparam \reg_file[26][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N18
cycloneive_lcell_comb \Mux55~2 (
// Equation(s):
// \Mux55~2_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[26][8]~q ))) # (!\prif.imemload_id [19] & (\reg_file[18][8]~q ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[18][8]~q ),
	.datac(\reg_file[26][8]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux55~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~2 .lut_mask = 16'hFA44;
defparam \Mux55~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N13
dffeas \reg_file[22][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][8] .is_wysiwyg = "true";
defparam \reg_file[22][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N12
cycloneive_lcell_comb \Mux55~3 (
// Equation(s):
// \Mux55~3_combout  = (\Mux55~2_combout  & ((\reg_file[30][8]~q ) # ((!\prif.imemload_id [18])))) # (!\Mux55~2_combout  & (((\reg_file[22][8]~q  & \prif.imemload_id [18]))))

	.dataa(\reg_file[30][8]~q ),
	.datab(\Mux55~2_combout ),
	.datac(\reg_file[22][8]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux55~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~3 .lut_mask = 16'hB8CC;
defparam \Mux55~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y26_N16
cycloneive_lcell_comb \Mux55~6 (
// Equation(s):
// \Mux55~6_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16]) # (\Mux55~3_combout )))) # (!\prif.imemload_id [17] & (\Mux55~5_combout  & (!\prif.imemload_id [16])))

	.dataa(prifimemload_id_17),
	.datab(\Mux55~5_combout ),
	.datac(prifimemload_id_16),
	.datad(\Mux55~3_combout ),
	.cin(gnd),
	.combout(\Mux55~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~6 .lut_mask = 16'hAEA4;
defparam \Mux55~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N8
cycloneive_lcell_comb \reg_file[2][8]~feeder (
// Equation(s):
// \reg_file[2][8]~feeder_combout  = \reg_file_nxt[31][8]~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][8]~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[2][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][8]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[2][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y26_N9
dffeas \reg_file[2][8] (
	.clk(!CLK),
	.d(\reg_file[2][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][8] .is_wysiwyg = "true";
defparam \reg_file[2][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N21
dffeas \reg_file[1][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][8] .is_wysiwyg = "true";
defparam \reg_file[1][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N11
dffeas \reg_file[3][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][8] .is_wysiwyg = "true";
defparam \reg_file[3][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N10
cycloneive_lcell_comb \Mux55~14 (
// Equation(s):
// \Mux55~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][8]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][8]~q ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[1][8]~q ),
	.datac(\reg_file[3][8]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux55~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~14 .lut_mask = 16'hE400;
defparam \Mux55~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N22
cycloneive_lcell_comb \Mux55~15 (
// Equation(s):
// \Mux55~15_combout  = (\Mux55~14_combout ) # ((!\prif.imemload_id [16] & (\prif.imemload_id [17] & \reg_file[2][8]~q )))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[2][8]~q ),
	.datad(\Mux55~14_combout ),
	.cin(gnd),
	.combout(\Mux55~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~15 .lut_mask = 16'hFF40;
defparam \Mux55~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y26_N23
dffeas \reg_file[6][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][8] .is_wysiwyg = "true";
defparam \reg_file[6][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N9
dffeas \reg_file[5][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][8] .is_wysiwyg = "true";
defparam \reg_file[5][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y26_N15
dffeas \reg_file[4][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][8] .is_wysiwyg = "true";
defparam \reg_file[4][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N14
cycloneive_lcell_comb \Mux55~12 (
// Equation(s):
// \Mux55~12_combout  = (\prif.imemload_id [16] & ((\reg_file[5][8]~q ) # ((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & (((\reg_file[4][8]~q  & !\prif.imemload_id [17]))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[5][8]~q ),
	.datac(\reg_file[4][8]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux55~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~12 .lut_mask = 16'hAAD8;
defparam \Mux55~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N18
cycloneive_lcell_comb \Mux55~13 (
// Equation(s):
// \Mux55~13_combout  = (\prif.imemload_id [17] & ((\Mux55~12_combout  & (\reg_file[7][8]~q )) # (!\Mux55~12_combout  & ((\reg_file[6][8]~q ))))) # (!\prif.imemload_id [17] & (((\Mux55~12_combout ))))

	.dataa(\reg_file[7][8]~q ),
	.datab(\reg_file[6][8]~q ),
	.datac(prifimemload_id_17),
	.datad(\Mux55~12_combout ),
	.cin(gnd),
	.combout(\Mux55~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~13 .lut_mask = 16'hAFC0;
defparam \Mux55~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N0
cycloneive_lcell_comb \Mux55~16 (
// Equation(s):
// \Mux55~16_combout  = (\prif.imemload_id [18] & (((\Mux55~13_combout ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\Mux55~15_combout  & ((!\prif.imemload_id [19]))))

	.dataa(\Mux55~15_combout ),
	.datab(\Mux55~13_combout ),
	.datac(prifimemload_id_18),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux55~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~16 .lut_mask = 16'hF0CA;
defparam \Mux55~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N23
dffeas \reg_file[8][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][8] .is_wysiwyg = "true";
defparam \reg_file[8][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N25
dffeas \reg_file[10][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][8] .is_wysiwyg = "true";
defparam \reg_file[10][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N22
cycloneive_lcell_comb \Mux55~10 (
// Equation(s):
// \Mux55~10_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\reg_file[10][8]~q )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & (\reg_file[8][8]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[8][8]~q ),
	.datad(\reg_file[10][8]~q ),
	.cin(gnd),
	.combout(\Mux55~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~10 .lut_mask = 16'hBA98;
defparam \Mux55~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N15
dffeas \reg_file[11][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][8] .is_wysiwyg = "true";
defparam \reg_file[11][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y33_N13
dffeas \reg_file[9][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][8] .is_wysiwyg = "true";
defparam \reg_file[9][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N12
cycloneive_lcell_comb \Mux55~11 (
// Equation(s):
// \Mux55~11_combout  = (\Mux55~10_combout  & ((\reg_file[11][8]~q ) # ((!\prif.imemload_id [16])))) # (!\Mux55~10_combout  & (((\reg_file[9][8]~q  & \prif.imemload_id [16]))))

	.dataa(\Mux55~10_combout ),
	.datab(\reg_file[11][8]~q ),
	.datac(\reg_file[9][8]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux55~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~11 .lut_mask = 16'hD8AA;
defparam \Mux55~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N2
cycloneive_lcell_comb \reg_file[15][8]~feeder (
// Equation(s):
// \reg_file[15][8]~feeder_combout  = \reg_file_nxt[31][8]~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][8]~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[15][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[15][8]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[15][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y27_N3
dffeas \reg_file[15][8] (
	.clk(!CLK),
	.d(\reg_file[15][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][8] .is_wysiwyg = "true";
defparam \reg_file[15][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y27_N29
dffeas \reg_file[14][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][8] .is_wysiwyg = "true";
defparam \reg_file[14][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N27
dffeas \reg_file[12][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][8] .is_wysiwyg = "true";
defparam \reg_file[12][8] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N5
dffeas \reg_file[13][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][8] .is_wysiwyg = "true";
defparam \reg_file[13][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N26
cycloneive_lcell_comb \Mux55~17 (
// Equation(s):
// \Mux55~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][8]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][8]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][8]~q ),
	.datad(\reg_file[13][8]~q ),
	.cin(gnd),
	.combout(\Mux55~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~17 .lut_mask = 16'hDC98;
defparam \Mux55~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N28
cycloneive_lcell_comb \Mux55~18 (
// Equation(s):
// \Mux55~18_combout  = (\prif.imemload_id [17] & ((\Mux55~17_combout  & (\reg_file[15][8]~q )) # (!\Mux55~17_combout  & ((\reg_file[14][8]~q ))))) # (!\prif.imemload_id [17] & (((\Mux55~17_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[15][8]~q ),
	.datac(\reg_file[14][8]~q ),
	.datad(\Mux55~17_combout ),
	.cin(gnd),
	.combout(\Mux55~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux55~18 .lut_mask = 16'hDDA0;
defparam \Mux55~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N10
cycloneive_lcell_comb \reg_file_nxt[31][7]~93 (
// Equation(s):
// \reg_file_nxt[31][7]~93_combout  = (\Mux157~1_combout  & (((\prif.regwrite_wb [0]) # (\prif.regwrite_wb [2])) # (!Equal8)))

	.dataa(Mux157),
	.datab(Equal8),
	.datac(prifregwrite_wb_0),
	.datad(prifregwrite_wb_2),
	.cin(gnd),
	.combout(\reg_file_nxt[31][7]~93_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][7]~93 .lut_mask = 16'hAAA2;
defparam \reg_file_nxt[31][7]~93 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y27_N13
dffeas \reg_file[19][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][7] .is_wysiwyg = "true";
defparam \reg_file[19][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y28_N31
dffeas \reg_file[27][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][7] .is_wysiwyg = "true";
defparam \reg_file[27][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N30
cycloneive_lcell_comb \Mux56~7 (
// Equation(s):
// \Mux56~7_combout  = (\prif.imemload_id [18] & (((\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\reg_file[27][7]~q ))) # (!\prif.imemload_id [19] & (\reg_file[19][7]~q ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[19][7]~q ),
	.datac(\reg_file[27][7]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux56~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~7 .lut_mask = 16'hFA44;
defparam \Mux56~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N24
cycloneive_lcell_comb \reg_file[23][7]~feeder (
// Equation(s):
// \reg_file[23][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][7]~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[23][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][7]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[23][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N25
dffeas \reg_file[23][7] (
	.clk(!CLK),
	.d(\reg_file[23][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][7] .is_wysiwyg = "true";
defparam \reg_file[23][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y27_N7
dffeas \reg_file[31][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][7] .is_wysiwyg = "true";
defparam \reg_file[31][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N0
cycloneive_lcell_comb \Mux56~8 (
// Equation(s):
// \Mux56~8_combout  = (\Mux56~7_combout  & (((\reg_file[31][7]~q )) # (!\prif.imemload_id [18]))) # (!\Mux56~7_combout  & (\prif.imemload_id [18] & (\reg_file[23][7]~q )))

	.dataa(\Mux56~7_combout ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[23][7]~q ),
	.datad(\reg_file[31][7]~q ),
	.cin(gnd),
	.combout(\Mux56~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~8 .lut_mask = 16'hEA62;
defparam \Mux56~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N12
cycloneive_lcell_comb \reg_file[29][7]~feeder (
// Equation(s):
// \reg_file[29][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][7]~93_combout ),
	.cin(gnd),
	.combout(\reg_file[29][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][7]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[29][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y32_N13
dffeas \reg_file[29][7] (
	.clk(!CLK),
	.d(\reg_file[29][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][7] .is_wysiwyg = "true";
defparam \reg_file[29][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y24_N12
cycloneive_lcell_comb \reg_file[21][7]~feeder (
// Equation(s):
// \reg_file[21][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][7]~93_combout ),
	.cin(gnd),
	.combout(\reg_file[21][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][7]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[21][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y24_N13
dffeas \reg_file[21][7] (
	.clk(!CLK),
	.d(\reg_file[21][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][7] .is_wysiwyg = "true";
defparam \reg_file[21][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N30
cycloneive_lcell_comb \reg_file[17][7]~feeder (
// Equation(s):
// \reg_file[17][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][7]~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[17][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[17][7]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[17][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y26_N31
dffeas \reg_file[17][7] (
	.clk(!CLK),
	.d(\reg_file[17][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][7] .is_wysiwyg = "true";
defparam \reg_file[17][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N31
dffeas \reg_file[25][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][7] .is_wysiwyg = "true";
defparam \reg_file[25][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N30
cycloneive_lcell_comb \Mux56~0 (
// Equation(s):
// \Mux56~0_combout  = (\prif.imemload_id [19] & (((\reg_file[25][7]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[17][7]~q  & ((!\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[17][7]~q ),
	.datac(\reg_file[25][7]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux56~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~0 .lut_mask = 16'hAAE4;
defparam \Mux56~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N2
cycloneive_lcell_comb \Mux56~1 (
// Equation(s):
// \Mux56~1_combout  = (\prif.imemload_id [18] & ((\Mux56~0_combout  & (\reg_file[29][7]~q )) # (!\Mux56~0_combout  & ((\reg_file[21][7]~q ))))) # (!\prif.imemload_id [18] & (((\Mux56~0_combout ))))

	.dataa(\reg_file[29][7]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[21][7]~q ),
	.datad(\Mux56~0_combout ),
	.cin(gnd),
	.combout(\Mux56~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~1 .lut_mask = 16'hBBC0;
defparam \Mux56~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N29
dffeas \reg_file[24][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][7] .is_wysiwyg = "true";
defparam \reg_file[24][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N28
cycloneive_lcell_comb \reg_file[20][7]~feeder (
// Equation(s):
// \reg_file[20][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][7]~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[20][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[20][7]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[20][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N29
dffeas \reg_file[20][7] (
	.clk(!CLK),
	.d(\reg_file[20][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][7] .is_wysiwyg = "true";
defparam \reg_file[20][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N16
cycloneive_lcell_comb \Mux56~4 (
// Equation(s):
// \Mux56~4_combout  = (\prif.imemload_id [18] & (((\reg_file[20][7]~q ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\reg_file[16][7]~q  & ((!\prif.imemload_id [19]))))

	.dataa(\reg_file[16][7]~q ),
	.datab(\reg_file[20][7]~q ),
	.datac(prifimemload_id_18),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux56~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~4 .lut_mask = 16'hF0CA;
defparam \Mux56~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N19
dffeas \reg_file[28][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][7] .is_wysiwyg = "true";
defparam \reg_file[28][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N0
cycloneive_lcell_comb \Mux56~5 (
// Equation(s):
// \Mux56~5_combout  = (\prif.imemload_id [19] & ((\Mux56~4_combout  & ((\reg_file[28][7]~q ))) # (!\Mux56~4_combout  & (\reg_file[24][7]~q )))) # (!\prif.imemload_id [19] & (((\Mux56~4_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[24][7]~q ),
	.datac(\Mux56~4_combout ),
	.datad(\reg_file[28][7]~q ),
	.cin(gnd),
	.combout(\Mux56~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~5 .lut_mask = 16'hF858;
defparam \Mux56~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N5
dffeas \reg_file[22][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][7] .is_wysiwyg = "true";
defparam \reg_file[22][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N4
cycloneive_lcell_comb \Mux56~2 (
// Equation(s):
// \Mux56~2_combout  = (\prif.imemload_id [18] & (((\reg_file[22][7]~q ) # (\prif.imemload_id [19])))) # (!\prif.imemload_id [18] & (\reg_file[18][7]~q  & ((!\prif.imemload_id [19]))))

	.dataa(\reg_file[18][7]~q ),
	.datab(prifimemload_id_18),
	.datac(\reg_file[22][7]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux56~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~2 .lut_mask = 16'hCCE2;
defparam \Mux56~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N1
dffeas \reg_file[26][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][7] .is_wysiwyg = "true";
defparam \reg_file[26][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N30
cycloneive_lcell_comb \reg_file[30][7]~feeder (
// Equation(s):
// \reg_file[30][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][7]~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[30][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[30][7]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[30][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N31
dffeas \reg_file[30][7] (
	.clk(!CLK),
	.d(\reg_file[30][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][7] .is_wysiwyg = "true";
defparam \reg_file[30][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N0
cycloneive_lcell_comb \Mux56~3 (
// Equation(s):
// \Mux56~3_combout  = (\prif.imemload_id [19] & ((\Mux56~2_combout  & ((\reg_file[30][7]~q ))) # (!\Mux56~2_combout  & (\reg_file[26][7]~q )))) # (!\prif.imemload_id [19] & (\Mux56~2_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux56~2_combout ),
	.datac(\reg_file[26][7]~q ),
	.datad(\reg_file[30][7]~q ),
	.cin(gnd),
	.combout(\Mux56~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~3 .lut_mask = 16'hEC64;
defparam \Mux56~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N24
cycloneive_lcell_comb \Mux56~6 (
// Equation(s):
// \Mux56~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux56~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & (\Mux56~5_combout )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux56~5_combout ),
	.datad(\Mux56~3_combout ),
	.cin(gnd),
	.combout(\Mux56~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~6 .lut_mask = 16'hBA98;
defparam \Mux56~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y28_N15
dffeas \reg_file[4][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][7] .is_wysiwyg = "true";
defparam \reg_file[4][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y28_N13
dffeas \reg_file[5][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][7] .is_wysiwyg = "true";
defparam \reg_file[5][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N12
cycloneive_lcell_comb \Mux56~10 (
// Equation(s):
// \Mux56~10_combout  = (\prif.imemload_id [17] & (((\prif.imemload_id [16])))) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[5][7]~q ))) # (!\prif.imemload_id [16] & (\reg_file[4][7]~q ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[4][7]~q ),
	.datac(\reg_file[5][7]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux56~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~10 .lut_mask = 16'hFA44;
defparam \Mux56~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N17
dffeas \reg_file[6][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][7] .is_wysiwyg = "true";
defparam \reg_file[6][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N11
dffeas \reg_file[7][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][7] .is_wysiwyg = "true";
defparam \reg_file[7][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N16
cycloneive_lcell_comb \Mux56~11 (
// Equation(s):
// \Mux56~11_combout  = (\prif.imemload_id [17] & ((\Mux56~10_combout  & ((\reg_file[7][7]~q ))) # (!\Mux56~10_combout  & (\reg_file[6][7]~q )))) # (!\prif.imemload_id [17] & (\Mux56~10_combout ))

	.dataa(prifimemload_id_17),
	.datab(\Mux56~10_combout ),
	.datac(\reg_file[6][7]~q ),
	.datad(\reg_file[7][7]~q ),
	.cin(gnd),
	.combout(\Mux56~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~11 .lut_mask = 16'hEC64;
defparam \Mux56~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y25_N31
dffeas \reg_file[12][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][7] .is_wysiwyg = "true";
defparam \reg_file[12][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y25_N29
dffeas \reg_file[13][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][7] .is_wysiwyg = "true";
defparam \reg_file[13][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N30
cycloneive_lcell_comb \Mux56~17 (
// Equation(s):
// \Mux56~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & ((\reg_file[13][7]~q ))) # (!\prif.imemload_id [16] & (\reg_file[12][7]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[12][7]~q ),
	.datad(\reg_file[13][7]~q ),
	.cin(gnd),
	.combout(\Mux56~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~17 .lut_mask = 16'hDC98;
defparam \Mux56~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N8
cycloneive_lcell_comb \reg_file[15][7]~feeder (
// Equation(s):
// \reg_file[15][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][7]~93_combout ),
	.cin(gnd),
	.combout(\reg_file[15][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[15][7]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[15][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y24_N9
dffeas \reg_file[15][7] (
	.clk(!CLK),
	.d(\reg_file[15][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][7] .is_wysiwyg = "true";
defparam \reg_file[15][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N20
cycloneive_lcell_comb \reg_file[14][7]~feeder (
// Equation(s):
// \reg_file[14][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][7]~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[14][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[14][7]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[14][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y26_N21
dffeas \reg_file[14][7] (
	.clk(!CLK),
	.d(\reg_file[14][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][7] .is_wysiwyg = "true";
defparam \reg_file[14][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N10
cycloneive_lcell_comb \Mux56~18 (
// Equation(s):
// \Mux56~18_combout  = (\Mux56~17_combout  & (((\reg_file[15][7]~q )) # (!\prif.imemload_id [17]))) # (!\Mux56~17_combout  & (\prif.imemload_id [17] & ((\reg_file[14][7]~q ))))

	.dataa(\Mux56~17_combout ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[15][7]~q ),
	.datad(\reg_file[14][7]~q ),
	.cin(gnd),
	.combout(\Mux56~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~18 .lut_mask = 16'hE6A2;
defparam \Mux56~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N28
cycloneive_lcell_comb \reg_file[2][7]~feeder (
// Equation(s):
// \reg_file[2][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][7]~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[2][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][7]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[2][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N29
dffeas \reg_file[2][7] (
	.clk(!CLK),
	.d(\reg_file[2][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][7] .is_wysiwyg = "true";
defparam \reg_file[2][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N21
dffeas \reg_file[1][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][7] .is_wysiwyg = "true";
defparam \reg_file[1][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X63_Y33_N11
dffeas \reg_file[3][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][7] .is_wysiwyg = "true";
defparam \reg_file[3][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N20
cycloneive_lcell_comb \Mux56~14 (
// Equation(s):
// \Mux56~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[3][7]~q ))) # (!\prif.imemload_id [17] & (\reg_file[1][7]~q ))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[1][7]~q ),
	.datad(\reg_file[3][7]~q ),
	.cin(gnd),
	.combout(\Mux56~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~14 .lut_mask = 16'hC840;
defparam \Mux56~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N26
cycloneive_lcell_comb \Mux56~15 (
// Equation(s):
// \Mux56~15_combout  = (\Mux56~14_combout ) # ((\prif.imemload_id [17] & (\reg_file[2][7]~q  & !\prif.imemload_id [16])))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[2][7]~q ),
	.datac(\Mux56~14_combout ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux56~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~15 .lut_mask = 16'hF0F8;
defparam \Mux56~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N0
cycloneive_lcell_comb \reg_file[11][7]~feeder (
// Equation(s):
// \reg_file[11][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][7]~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[11][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[11][7]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[11][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y35_N1
dffeas \reg_file[11][7] (
	.clk(!CLK),
	.d(\reg_file[11][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][7] .is_wysiwyg = "true";
defparam \reg_file[11][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N7
dffeas \reg_file[8][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][7] .is_wysiwyg = "true";
defparam \reg_file[8][7] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N1
dffeas \reg_file[10][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][7] .is_wysiwyg = "true";
defparam \reg_file[10][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N6
cycloneive_lcell_comb \Mux56~12 (
// Equation(s):
// \Mux56~12_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\reg_file[10][7]~q )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & (\reg_file[8][7]~q )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[8][7]~q ),
	.datad(\reg_file[10][7]~q ),
	.cin(gnd),
	.combout(\Mux56~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~12 .lut_mask = 16'hBA98;
defparam \Mux56~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N10
cycloneive_lcell_comb \Mux56~13 (
// Equation(s):
// \Mux56~13_combout  = (\Mux56~12_combout  & (((\reg_file[11][7]~q ) # (!\prif.imemload_id [16])))) # (!\Mux56~12_combout  & (\reg_file[9][7]~q  & ((\prif.imemload_id [16]))))

	.dataa(\reg_file[9][7]~q ),
	.datab(\reg_file[11][7]~q ),
	.datac(\Mux56~12_combout ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux56~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~13 .lut_mask = 16'hCAF0;
defparam \Mux56~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y35_N16
cycloneive_lcell_comb \Mux56~16 (
// Equation(s):
// \Mux56~16_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & ((\Mux56~13_combout ))) # (!\prif.imemload_id [19] & (\Mux56~15_combout ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\Mux56~15_combout ),
	.datad(\Mux56~13_combout ),
	.cin(gnd),
	.combout(\Mux56~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux56~16 .lut_mask = 16'hDC98;
defparam \Mux56~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N0
cycloneive_lcell_comb \reg_file_nxt[31][22]~94 (
// Equation(s):
// \reg_file_nxt[31][22]~94_combout  = (\Mux142~1_combout  & (((\prif.regwrite_wb [2]) # (\prif.regwrite_wb [0])) # (!Equal8)))

	.dataa(Equal8),
	.datab(prifregwrite_wb_2),
	.datac(Mux142),
	.datad(prifregwrite_wb_0),
	.cin(gnd),
	.combout(\reg_file_nxt[31][22]~94_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][22]~94 .lut_mask = 16'hF0D0;
defparam \reg_file_nxt[31][22]~94 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N6
cycloneive_lcell_comb \reg_file[29][22]~feeder (
// Equation(s):
// \reg_file[29][22]~feeder_combout  = \reg_file_nxt[31][22]~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][22]~94_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][22]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N7
dffeas \reg_file[29][22] (
	.clk(!CLK),
	.d(\reg_file[29][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][22] .is_wysiwyg = "true";
defparam \reg_file[29][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N15
dffeas \reg_file[25][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][22] .is_wysiwyg = "true";
defparam \reg_file[25][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y30_N17
dffeas \reg_file[17][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][22] .is_wysiwyg = "true";
defparam \reg_file[17][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N1
dffeas \reg_file[21][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][22] .is_wysiwyg = "true";
defparam \reg_file[21][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N0
cycloneive_lcell_comb \Mux41~0 (
// Equation(s):
// \Mux41~0_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[21][22]~q ))) # (!\prif.imemload_id [18] & (\reg_file[17][22]~q ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[17][22]~q ),
	.datac(\reg_file[21][22]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux41~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~0 .lut_mask = 16'hFA44;
defparam \Mux41~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N14
cycloneive_lcell_comb \Mux41~1 (
// Equation(s):
// \Mux41~1_combout  = (\prif.imemload_id [19] & ((\Mux41~0_combout  & (\reg_file[29][22]~q )) # (!\Mux41~0_combout  & ((\reg_file[25][22]~q ))))) # (!\prif.imemload_id [19] & (((\Mux41~0_combout ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[29][22]~q ),
	.datac(\reg_file[25][22]~q ),
	.datad(\Mux41~0_combout ),
	.cin(gnd),
	.combout(\Mux41~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~1 .lut_mask = 16'hDDA0;
defparam \Mux41~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N12
cycloneive_lcell_comb \reg_file[27][22]~feeder (
// Equation(s):
// \reg_file[27][22]~feeder_combout  = \reg_file_nxt[31][22]~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][22]~94_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[27][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[27][22]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[27][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N13
dffeas \reg_file[27][22] (
	.clk(!CLK),
	.d(\reg_file[27][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][22] .is_wysiwyg = "true";
defparam \reg_file[27][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N1
dffeas \reg_file[31][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][22] .is_wysiwyg = "true";
defparam \reg_file[31][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y29_N19
dffeas \reg_file[23][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][22] .is_wysiwyg = "true";
defparam \reg_file[23][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y29_N31
dffeas \reg_file[19][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][22] .is_wysiwyg = "true";
defparam \reg_file[19][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N18
cycloneive_lcell_comb \Mux41~7 (
// Equation(s):
// \Mux41~7_combout  = (\prif.imemload_id [18] & ((\prif.imemload_id [19]) # ((\reg_file[23][22]~q )))) # (!\prif.imemload_id [18] & (!\prif.imemload_id [19] & ((\reg_file[19][22]~q ))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[23][22]~q ),
	.datad(\reg_file[19][22]~q ),
	.cin(gnd),
	.combout(\Mux41~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~7 .lut_mask = 16'hB9A8;
defparam \Mux41~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N0
cycloneive_lcell_comb \Mux41~8 (
// Equation(s):
// \Mux41~8_combout  = (\prif.imemload_id [19] & ((\Mux41~7_combout  & ((\reg_file[31][22]~q ))) # (!\Mux41~7_combout  & (\reg_file[27][22]~q )))) # (!\prif.imemload_id [19] & (((\Mux41~7_combout ))))

	.dataa(\reg_file[27][22]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[31][22]~q ),
	.datad(\Mux41~7_combout ),
	.cin(gnd),
	.combout(\Mux41~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~8 .lut_mask = 16'hF388;
defparam \Mux41~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N15
dffeas \reg_file[28][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][22] .is_wysiwyg = "true";
defparam \reg_file[28][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N13
dffeas \reg_file[20][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][22] .is_wysiwyg = "true";
defparam \reg_file[20][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y33_N17
dffeas \reg_file[24][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][22] .is_wysiwyg = "true";
defparam \reg_file[24][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N16
cycloneive_lcell_comb \Mux41~4 (
// Equation(s):
// \Mux41~4_combout  = (\prif.imemload_id [19] & (((\reg_file[24][22]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[16][22]~q  & ((!\prif.imemload_id [18]))))

	.dataa(\reg_file[16][22]~q ),
	.datab(prifimemload_id_19),
	.datac(\reg_file[24][22]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux41~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~4 .lut_mask = 16'hCCE2;
defparam \Mux41~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N12
cycloneive_lcell_comb \Mux41~5 (
// Equation(s):
// \Mux41~5_combout  = (\prif.imemload_id [18] & ((\Mux41~4_combout  & (\reg_file[28][22]~q )) # (!\Mux41~4_combout  & ((\reg_file[20][22]~q ))))) # (!\prif.imemload_id [18] & (((\Mux41~4_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[28][22]~q ),
	.datac(\reg_file[20][22]~q ),
	.datad(\Mux41~4_combout ),
	.cin(gnd),
	.combout(\Mux41~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~5 .lut_mask = 16'hDDA0;
defparam \Mux41~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N30
cycloneive_lcell_comb \reg_file[22][22]~feeder (
// Equation(s):
// \reg_file[22][22]~feeder_combout  = \reg_file_nxt[31][22]~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][22]~94_combout ),
	.cin(gnd),
	.combout(\reg_file[22][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][22]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[22][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N31
dffeas \reg_file[22][22] (
	.clk(!CLK),
	.d(\reg_file[22][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][22] .is_wysiwyg = "true";
defparam \reg_file[22][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y28_N7
dffeas \reg_file[30][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][22] .is_wysiwyg = "true";
defparam \reg_file[30][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y30_N27
dffeas \reg_file[18][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][22] .is_wysiwyg = "true";
defparam \reg_file[18][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y30_N17
dffeas \reg_file[26][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][22] .is_wysiwyg = "true";
defparam \reg_file[26][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N16
cycloneive_lcell_comb \Mux41~2 (
// Equation(s):
// \Mux41~2_combout  = (\prif.imemload_id [19] & (((\reg_file[26][22]~q ) # (\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & (\reg_file[18][22]~q  & ((!\prif.imemload_id [18]))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[18][22]~q ),
	.datac(\reg_file[26][22]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux41~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~2 .lut_mask = 16'hAAE4;
defparam \Mux41~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N6
cycloneive_lcell_comb \Mux41~3 (
// Equation(s):
// \Mux41~3_combout  = (\prif.imemload_id [18] & ((\Mux41~2_combout  & ((\reg_file[30][22]~q ))) # (!\Mux41~2_combout  & (\reg_file[22][22]~q )))) # (!\prif.imemload_id [18] & (((\Mux41~2_combout ))))

	.dataa(prifimemload_id_18),
	.datab(\reg_file[22][22]~q ),
	.datac(\reg_file[30][22]~q ),
	.datad(\Mux41~2_combout ),
	.cin(gnd),
	.combout(\Mux41~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~3 .lut_mask = 16'hF588;
defparam \Mux41~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N24
cycloneive_lcell_comb \Mux41~6 (
// Equation(s):
// \Mux41~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux41~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & (\Mux41~5_combout )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux41~5_combout ),
	.datad(\Mux41~3_combout ),
	.cin(gnd),
	.combout(\Mux41~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~6 .lut_mask = 16'hBA98;
defparam \Mux41~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N9
dffeas \reg_file[13][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][22] .is_wysiwyg = "true";
defparam \reg_file[13][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y32_N23
dffeas \reg_file[12][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][22] .is_wysiwyg = "true";
defparam \reg_file[12][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N22
cycloneive_lcell_comb \Mux41~17 (
// Equation(s):
// \Mux41~17_combout  = (\prif.imemload_id [16] & ((\reg_file[13][22]~q ) # ((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & (((\reg_file[12][22]~q  & !\prif.imemload_id [17]))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[13][22]~q ),
	.datac(\reg_file[12][22]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux41~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~17 .lut_mask = 16'hAAD8;
defparam \Mux41~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N11
dffeas \reg_file[14][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][22] .is_wysiwyg = "true";
defparam \reg_file[14][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y31_N1
dffeas \reg_file[15][22] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][22]~94_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][22] .is_wysiwyg = "true";
defparam \reg_file[15][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N10
cycloneive_lcell_comb \Mux41~18 (
// Equation(s):
// \Mux41~18_combout  = (\prif.imemload_id [17] & ((\Mux41~17_combout  & ((\reg_file[15][22]~q ))) # (!\Mux41~17_combout  & (\reg_file[14][22]~q )))) # (!\prif.imemload_id [17] & (\Mux41~17_combout ))

	.dataa(prifimemload_id_17),
	.datab(\Mux41~17_combout ),
	.datac(\reg_file[14][22]~q ),
	.datad(\reg_file[15][22]~q ),
	.cin(gnd),
	.combout(\Mux41~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~18 .lut_mask = 16'hEC64;
defparam \Mux41~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N19
dffeas \reg_file[11][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][22] .is_wysiwyg = "true";
defparam \reg_file[11][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X68_Y35_N5
dffeas \reg_file[9][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][22] .is_wysiwyg = "true";
defparam \reg_file[9][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N7
dffeas \reg_file[8][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][22] .is_wysiwyg = "true";
defparam \reg_file[8][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y35_N17
dffeas \reg_file[10][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][22] .is_wysiwyg = "true";
defparam \reg_file[10][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N6
cycloneive_lcell_comb \Mux41~10 (
// Equation(s):
// \Mux41~10_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][22]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][22]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[8][22]~q ),
	.datad(\reg_file[10][22]~q ),
	.cin(gnd),
	.combout(\Mux41~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~10 .lut_mask = 16'hDC98;
defparam \Mux41~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N4
cycloneive_lcell_comb \Mux41~11 (
// Equation(s):
// \Mux41~11_combout  = (\prif.imemload_id [16] & ((\Mux41~10_combout  & (\reg_file[11][22]~q )) # (!\Mux41~10_combout  & ((\reg_file[9][22]~q ))))) # (!\prif.imemload_id [16] & (((\Mux41~10_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[11][22]~q ),
	.datac(\reg_file[9][22]~q ),
	.datad(\Mux41~10_combout ),
	.cin(gnd),
	.combout(\Mux41~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~11 .lut_mask = 16'hDDA0;
defparam \Mux41~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y32_N19
dffeas \reg_file[3][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][22] .is_wysiwyg = "true";
defparam \reg_file[3][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y32_N13
dffeas \reg_file[1][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][22] .is_wysiwyg = "true";
defparam \reg_file[1][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N12
cycloneive_lcell_comb \Mux41~14 (
// Equation(s):
// \Mux41~14_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17] & (\reg_file[3][22]~q )) # (!\prif.imemload_id [17] & ((\reg_file[1][22]~q )))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[3][22]~q ),
	.datac(\reg_file[1][22]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux41~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~14 .lut_mask = 16'hD800;
defparam \Mux41~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N11
dffeas \reg_file[2][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][22] .is_wysiwyg = "true";
defparam \reg_file[2][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N10
cycloneive_lcell_comb \Mux41~15 (
// Equation(s):
// \Mux41~15_combout  = (\Mux41~14_combout ) # ((\prif.imemload_id [17] & (\reg_file[2][22]~q  & !\prif.imemload_id [16])))

	.dataa(prifimemload_id_17),
	.datab(\Mux41~14_combout ),
	.datac(\reg_file[2][22]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux41~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~15 .lut_mask = 16'hCCEC;
defparam \Mux41~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N28
cycloneive_lcell_comb \reg_file[7][22]~feeder (
// Equation(s):
// \reg_file[7][22]~feeder_combout  = \reg_file_nxt[31][22]~94_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][22]~94_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[7][22]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[7][22]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[7][22]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N29
dffeas \reg_file[7][22] (
	.clk(!CLK),
	.d(\reg_file[7][22]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][22] .is_wysiwyg = "true";
defparam \reg_file[7][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N9
dffeas \reg_file[5][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][22] .is_wysiwyg = "true";
defparam \reg_file[5][22] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N31
dffeas \reg_file[4][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][22] .is_wysiwyg = "true";
defparam \reg_file[4][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N30
cycloneive_lcell_comb \Mux41~12 (
// Equation(s):
// \Mux41~12_combout  = (\prif.imemload_id [16] & ((\reg_file[5][22]~q ) # ((\prif.imemload_id [17])))) # (!\prif.imemload_id [16] & (((\reg_file[4][22]~q  & !\prif.imemload_id [17]))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[5][22]~q ),
	.datac(\reg_file[4][22]~q ),
	.datad(prifimemload_id_17),
	.cin(gnd),
	.combout(\Mux41~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~12 .lut_mask = 16'hAAD8;
defparam \Mux41~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y30_N17
dffeas \reg_file[6][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][22] .is_wysiwyg = "true";
defparam \reg_file[6][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N18
cycloneive_lcell_comb \Mux41~13 (
// Equation(s):
// \Mux41~13_combout  = (\prif.imemload_id [17] & ((\Mux41~12_combout  & (\reg_file[7][22]~q )) # (!\Mux41~12_combout  & ((\reg_file[6][22]~q ))))) # (!\prif.imemload_id [17] & (((\Mux41~12_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[7][22]~q ),
	.datac(\Mux41~12_combout ),
	.datad(\reg_file[6][22]~q ),
	.cin(gnd),
	.combout(\Mux41~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~13 .lut_mask = 16'hDAD0;
defparam \Mux41~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N16
cycloneive_lcell_comb \Mux41~16 (
// Equation(s):
// \Mux41~16_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\Mux41~13_combout ))) # (!\prif.imemload_id [18] & (\Mux41~15_combout ))))

	.dataa(\Mux41~15_combout ),
	.datab(prifimemload_id_19),
	.datac(prifimemload_id_18),
	.datad(\Mux41~13_combout ),
	.cin(gnd),
	.combout(\Mux41~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux41~16 .lut_mask = 16'hF2C2;
defparam \Mux41~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N18
cycloneive_lcell_comb \reg_file_nxt[31][25]~95 (
// Equation(s):
// \reg_file_nxt[31][25]~95_combout  = (\Mux139~1_combout  & ((\prif.regwrite_wb [2]) # ((\prif.regwrite_wb [0]) # (!Equal8))))

	.dataa(prifregwrite_wb_2),
	.datab(prifregwrite_wb_0),
	.datac(Mux139),
	.datad(Equal8),
	.cin(gnd),
	.combout(\reg_file_nxt[31][25]~95_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file_nxt[31][25]~95 .lut_mask = 16'hE0F0;
defparam \reg_file_nxt[31][25]~95 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N4
cycloneive_lcell_comb \reg_file[23][25]~feeder (
// Equation(s):
// \reg_file[23][25]~feeder_combout  = \reg_file_nxt[31][25]~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][25]~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[23][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[23][25]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[23][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N5
dffeas \reg_file[23][25] (
	.clk(!CLK),
	.d(\reg_file[23][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~30_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[23][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[23][25] .is_wysiwyg = "true";
defparam \reg_file[23][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y26_N5
dffeas \reg_file[27][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~31_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[27][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[27][25] .is_wysiwyg = "true";
defparam \reg_file[27][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y27_N21
dffeas \reg_file[19][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][25] .is_wysiwyg = "true";
defparam \reg_file[19][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N4
cycloneive_lcell_comb \Mux38~7 (
// Equation(s):
// \Mux38~7_combout  = (\prif.imemload_id [18] & (\prif.imemload_id [19])) # (!\prif.imemload_id [18] & ((\prif.imemload_id [19] & (\reg_file[27][25]~q )) # (!\prif.imemload_id [19] & ((\reg_file[19][25]~q )))))

	.dataa(prifimemload_id_18),
	.datab(prifimemload_id_19),
	.datac(\reg_file[27][25]~q ),
	.datad(\reg_file[19][25]~q ),
	.cin(gnd),
	.combout(\Mux38~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~7 .lut_mask = 16'hD9C8;
defparam \Mux38~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y26_N15
dffeas \reg_file[31][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~33_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[31][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[31][25] .is_wysiwyg = "true";
defparam \reg_file[31][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N14
cycloneive_lcell_comb \Mux38~8 (
// Equation(s):
// \Mux38~8_combout  = (\Mux38~7_combout  & (((\reg_file[31][25]~q ) # (!\prif.imemload_id [18])))) # (!\Mux38~7_combout  & (\reg_file[23][25]~q  & ((\prif.imemload_id [18]))))

	.dataa(\reg_file[23][25]~q ),
	.datab(\Mux38~7_combout ),
	.datac(\reg_file[31][25]~q ),
	.datad(prifimemload_id_18),
	.cin(gnd),
	.combout(\Mux38~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~8 .lut_mask = 16'hE2CC;
defparam \Mux38~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N3
dffeas \reg_file[25][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][25] .is_wysiwyg = "true";
defparam \reg_file[25][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N2
cycloneive_lcell_comb \reg_file[17][25]~feeder (
// Equation(s):
// \reg_file[17][25]~feeder_combout  = \reg_file_nxt[31][25]~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][25]~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[17][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[17][25]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[17][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y26_N3
dffeas \reg_file[17][25] (
	.clk(!CLK),
	.d(\reg_file[17][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][25] .is_wysiwyg = "true";
defparam \reg_file[17][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N2
cycloneive_lcell_comb \Mux38~0 (
// Equation(s):
// \Mux38~0_combout  = (\prif.imemload_id [19] & ((\prif.imemload_id [18]) # ((\reg_file[25][25]~q )))) # (!\prif.imemload_id [19] & (!\prif.imemload_id [18] & ((\reg_file[17][25]~q ))))

	.dataa(prifimemload_id_19),
	.datab(prifimemload_id_18),
	.datac(\reg_file[25][25]~q ),
	.datad(\reg_file[17][25]~q ),
	.cin(gnd),
	.combout(\Mux38~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~0 .lut_mask = 16'hB9A8;
defparam \Mux38~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y26_N27
dffeas \reg_file[21][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][25] .is_wysiwyg = "true";
defparam \reg_file[21][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N26
cycloneive_lcell_comb \reg_file[29][25]~feeder (
// Equation(s):
// \reg_file[29][25]~feeder_combout  = \reg_file_nxt[31][25]~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][25]~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[29][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[29][25]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[29][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y29_N27
dffeas \reg_file[29][25] (
	.clk(!CLK),
	.d(\reg_file[29][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~19_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[29][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[29][25] .is_wysiwyg = "true";
defparam \reg_file[29][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N26
cycloneive_lcell_comb \Mux38~1 (
// Equation(s):
// \Mux38~1_combout  = (\prif.imemload_id [18] & ((\Mux38~0_combout  & ((\reg_file[29][25]~q ))) # (!\Mux38~0_combout  & (\reg_file[21][25]~q )))) # (!\prif.imemload_id [18] & (\Mux38~0_combout ))

	.dataa(prifimemload_id_18),
	.datab(\Mux38~0_combout ),
	.datac(\reg_file[21][25]~q ),
	.datad(\reg_file[29][25]~q ),
	.cin(gnd),
	.combout(\Mux38~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~1 .lut_mask = 16'hEC64;
defparam \Mux38~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N25
dffeas \reg_file[28][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][25] .is_wysiwyg = "true";
defparam \reg_file[28][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y34_N11
dffeas \reg_file[24][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][25] .is_wysiwyg = "true";
defparam \reg_file[24][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N10
cycloneive_lcell_comb \Mux38~5 (
// Equation(s):
// \Mux38~5_combout  = (\Mux38~4_combout  & ((\reg_file[28][25]~q ) # ((!\prif.imemload_id [19])))) # (!\Mux38~4_combout  & (((\reg_file[24][25]~q  & \prif.imemload_id [19]))))

	.dataa(\Mux38~4_combout ),
	.datab(\reg_file[28][25]~q ),
	.datac(\reg_file[24][25]~q ),
	.datad(prifimemload_id_19),
	.cin(gnd),
	.combout(\Mux38~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~5 .lut_mask = 16'hD8AA;
defparam \Mux38~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N20
cycloneive_lcell_comb \reg_file[18][25]~feeder (
// Equation(s):
// \reg_file[18][25]~feeder_combout  = \reg_file_nxt[31][25]~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][25]~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[18][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[18][25]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[18][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N21
dffeas \reg_file[18][25] (
	.clk(!CLK),
	.d(\reg_file[18][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][25] .is_wysiwyg = "true";
defparam \reg_file[18][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N16
cycloneive_lcell_comb \reg_file[22][25]~feeder (
// Equation(s):
// \reg_file[22][25]~feeder_combout  = \reg_file_nxt[31][25]~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][25]~95_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[22][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][25]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[22][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y30_N17
dffeas \reg_file[22][25] (
	.clk(!CLK),
	.d(\reg_file[22][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][25] .is_wysiwyg = "true";
defparam \reg_file[22][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N2
cycloneive_lcell_comb \Mux38~2 (
// Equation(s):
// \Mux38~2_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18])))) # (!\prif.imemload_id [19] & ((\prif.imemload_id [18] & ((\reg_file[22][25]~q ))) # (!\prif.imemload_id [18] & (\reg_file[18][25]~q ))))

	.dataa(prifimemload_id_19),
	.datab(\reg_file[18][25]~q ),
	.datac(prifimemload_id_18),
	.datad(\reg_file[22][25]~q ),
	.cin(gnd),
	.combout(\Mux38~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~2 .lut_mask = 16'hF4A4;
defparam \Mux38~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y30_N17
dffeas \reg_file[30][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][25] .is_wysiwyg = "true";
defparam \reg_file[30][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N6
cycloneive_lcell_comb \reg_file[26][25]~feeder (
// Equation(s):
// \reg_file[26][25]~feeder_combout  = \reg_file_nxt[31][25]~95_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][25]~95_combout ),
	.cin(gnd),
	.combout(\reg_file[26][25]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[26][25]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[26][25]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N7
dffeas \reg_file[26][25] (
	.clk(!CLK),
	.d(\reg_file[26][25]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][25] .is_wysiwyg = "true";
defparam \reg_file[26][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N16
cycloneive_lcell_comb \Mux38~3 (
// Equation(s):
// \Mux38~3_combout  = (\prif.imemload_id [19] & ((\Mux38~2_combout  & (\reg_file[30][25]~q )) # (!\Mux38~2_combout  & ((\reg_file[26][25]~q ))))) # (!\prif.imemload_id [19] & (\Mux38~2_combout ))

	.dataa(prifimemload_id_19),
	.datab(\Mux38~2_combout ),
	.datac(\reg_file[30][25]~q ),
	.datad(\reg_file[26][25]~q ),
	.cin(gnd),
	.combout(\Mux38~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~3 .lut_mask = 16'hE6C4;
defparam \Mux38~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y30_N16
cycloneive_lcell_comb \Mux38~6 (
// Equation(s):
// \Mux38~6_combout  = (\prif.imemload_id [17] & ((\prif.imemload_id [16]) # ((\Mux38~3_combout )))) # (!\prif.imemload_id [17] & (!\prif.imemload_id [16] & (\Mux38~5_combout )))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\Mux38~5_combout ),
	.datad(\Mux38~3_combout ),
	.cin(gnd),
	.combout(\Mux38~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~6 .lut_mask = 16'hBA98;
defparam \Mux38~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y29_N19
dffeas \reg_file[15][25] (
	.clk(!CLK),
	.d(\reg_file_nxt[31][25]~95_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~41_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[15][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[15][25] .is_wysiwyg = "true";
defparam \reg_file[15][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y26_N13
dffeas \reg_file[14][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~38_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[14][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[14][25] .is_wysiwyg = "true";
defparam \reg_file[14][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N17
dffeas \reg_file[13][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~39_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[13][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[13][25] .is_wysiwyg = "true";
defparam \reg_file[13][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y26_N19
dffeas \reg_file[12][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][25] .is_wysiwyg = "true";
defparam \reg_file[12][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N16
cycloneive_lcell_comb \Mux38~17 (
// Equation(s):
// \Mux38~17_combout  = (\prif.imemload_id [17] & (\prif.imemload_id [16])) # (!\prif.imemload_id [17] & ((\prif.imemload_id [16] & (\reg_file[13][25]~q )) # (!\prif.imemload_id [16] & ((\reg_file[12][25]~q )))))

	.dataa(prifimemload_id_17),
	.datab(prifimemload_id_16),
	.datac(\reg_file[13][25]~q ),
	.datad(\reg_file[12][25]~q ),
	.cin(gnd),
	.combout(\Mux38~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~17 .lut_mask = 16'hD9C8;
defparam \Mux38~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N12
cycloneive_lcell_comb \Mux38~18 (
// Equation(s):
// \Mux38~18_combout  = (\prif.imemload_id [17] & ((\Mux38~17_combout  & (\reg_file[15][25]~q )) # (!\Mux38~17_combout  & ((\reg_file[14][25]~q ))))) # (!\prif.imemload_id [17] & (((\Mux38~17_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[15][25]~q ),
	.datac(\reg_file[14][25]~q ),
	.datad(\Mux38~17_combout ),
	.cin(gnd),
	.combout(\Mux38~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~18 .lut_mask = 16'hDDA0;
defparam \Mux38~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y34_N9
dffeas \reg_file[2][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][25] .is_wysiwyg = "true";
defparam \reg_file[2][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N0
cycloneive_lcell_comb \Mux38~15 (
// Equation(s):
// \Mux38~15_combout  = (\Mux38~14_combout ) # ((\prif.imemload_id [17] & (\reg_file[2][25]~q  & !\prif.imemload_id [16])))

	.dataa(\Mux38~14_combout ),
	.datab(prifimemload_id_17),
	.datac(\reg_file[2][25]~q ),
	.datad(prifimemload_id_16),
	.cin(gnd),
	.combout(\Mux38~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~15 .lut_mask = 16'hAAEA;
defparam \Mux38~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y25_N25
dffeas \reg_file[9][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][25] .is_wysiwyg = "true";
defparam \reg_file[9][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y25_N27
dffeas \reg_file[11][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][25] .is_wysiwyg = "true";
defparam \reg_file[11][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N7
dffeas \reg_file[8][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][25] .is_wysiwyg = "true";
defparam \reg_file[8][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X70_Y25_N29
dffeas \reg_file[10][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][25] .is_wysiwyg = "true";
defparam \reg_file[10][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N6
cycloneive_lcell_comb \Mux38~12 (
// Equation(s):
// \Mux38~12_combout  = (\prif.imemload_id [16] & (\prif.imemload_id [17])) # (!\prif.imemload_id [16] & ((\prif.imemload_id [17] & ((\reg_file[10][25]~q ))) # (!\prif.imemload_id [17] & (\reg_file[8][25]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[8][25]~q ),
	.datad(\reg_file[10][25]~q ),
	.cin(gnd),
	.combout(\Mux38~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~12 .lut_mask = 16'hDC98;
defparam \Mux38~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N26
cycloneive_lcell_comb \Mux38~13 (
// Equation(s):
// \Mux38~13_combout  = (\prif.imemload_id [16] & ((\Mux38~12_combout  & ((\reg_file[11][25]~q ))) # (!\Mux38~12_combout  & (\reg_file[9][25]~q )))) # (!\prif.imemload_id [16] & (((\Mux38~12_combout ))))

	.dataa(prifimemload_id_16),
	.datab(\reg_file[9][25]~q ),
	.datac(\reg_file[11][25]~q ),
	.datad(\Mux38~12_combout ),
	.cin(gnd),
	.combout(\Mux38~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~13 .lut_mask = 16'hF588;
defparam \Mux38~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N18
cycloneive_lcell_comb \Mux38~16 (
// Equation(s):
// \Mux38~16_combout  = (\prif.imemload_id [19] & (((\prif.imemload_id [18]) # (\Mux38~13_combout )))) # (!\prif.imemload_id [19] & (\Mux38~15_combout  & (!\prif.imemload_id [18])))

	.dataa(prifimemload_id_19),
	.datab(\Mux38~15_combout ),
	.datac(prifimemload_id_18),
	.datad(\Mux38~13_combout ),
	.cin(gnd),
	.combout(\Mux38~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~16 .lut_mask = 16'hAEA4;
defparam \Mux38~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N3
dffeas \reg_file[7][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][25] .is_wysiwyg = "true";
defparam \reg_file[7][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X72_Y28_N21
dffeas \reg_file[6][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][25] .is_wysiwyg = "true";
defparam \reg_file[6][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N25
dffeas \reg_file[5][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][25] .is_wysiwyg = "true";
defparam \reg_file[5][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N7
dffeas \reg_file[4][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][25] .is_wysiwyg = "true";
defparam \reg_file[4][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N24
cycloneive_lcell_comb \Mux38~10 (
// Equation(s):
// \Mux38~10_combout  = (\prif.imemload_id [16] & ((\prif.imemload_id [17]) # ((\reg_file[5][25]~q )))) # (!\prif.imemload_id [16] & (!\prif.imemload_id [17] & ((\reg_file[4][25]~q ))))

	.dataa(prifimemload_id_16),
	.datab(prifimemload_id_17),
	.datac(\reg_file[5][25]~q ),
	.datad(\reg_file[4][25]~q ),
	.cin(gnd),
	.combout(\Mux38~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~10 .lut_mask = 16'hB9A8;
defparam \Mux38~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N20
cycloneive_lcell_comb \Mux38~11 (
// Equation(s):
// \Mux38~11_combout  = (\prif.imemload_id [17] & ((\Mux38~10_combout  & (\reg_file[7][25]~q )) # (!\Mux38~10_combout  & ((\reg_file[6][25]~q ))))) # (!\prif.imemload_id [17] & (((\Mux38~10_combout ))))

	.dataa(prifimemload_id_17),
	.datab(\reg_file[7][25]~q ),
	.datac(\reg_file[6][25]~q ),
	.datad(\Mux38~10_combout ),
	.cin(gnd),
	.combout(\Mux38~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux38~11 .lut_mask = 16'hDDA0;
defparam \Mux38~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N2
cycloneive_lcell_comb \Mux29~0 (
// Equation(s):
// \Mux29~0_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][2]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][2]~q )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[25][2]~q ),
	.datad(\reg_file[17][2]~q ),
	.cin(gnd),
	.combout(\Mux29~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~0 .lut_mask = 16'hD9C8;
defparam \Mux29~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y24_N6
cycloneive_lcell_comb \Mux29~1 (
// Equation(s):
// \Mux29~1_combout  = (\prif.imemload_id [23] & ((\Mux29~0_combout  & (\reg_file[29][2]~q )) # (!\Mux29~0_combout  & ((\reg_file[21][2]~q ))))) # (!\prif.imemload_id [23] & (((\Mux29~0_combout ))))

	.dataa(\reg_file[29][2]~q ),
	.datab(\reg_file[21][2]~q ),
	.datac(prifimemload_id_23),
	.datad(\Mux29~0_combout ),
	.cin(gnd),
	.combout(\Mux29~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~1 .lut_mask = 16'hAFC0;
defparam \Mux29~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N20
cycloneive_lcell_comb \Mux29~7 (
// Equation(s):
// \Mux29~7_combout  = (\prif.imemload_id [24] & ((\reg_file[27][2]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[19][2]~q  & !\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[27][2]~q ),
	.datac(\reg_file[19][2]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux29~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~7 .lut_mask = 16'hAAD8;
defparam \Mux29~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N26
cycloneive_lcell_comb \Mux29~8 (
// Equation(s):
// \Mux29~8_combout  = (\prif.imemload_id [23] & ((\Mux29~7_combout  & ((\reg_file[31][2]~q ))) # (!\Mux29~7_combout  & (\reg_file[23][2]~q )))) # (!\prif.imemload_id [23] & (((\Mux29~7_combout ))))

	.dataa(\reg_file[23][2]~q ),
	.datab(\reg_file[31][2]~q ),
	.datac(prifimemload_id_23),
	.datad(\Mux29~7_combout ),
	.cin(gnd),
	.combout(\Mux29~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~8 .lut_mask = 16'hCFA0;
defparam \Mux29~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N23
dffeas \reg_file[28][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][2] .is_wysiwyg = "true";
defparam \reg_file[28][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N22
cycloneive_lcell_comb \Mux29~5 (
// Equation(s):
// \Mux29~5_combout  = (\Mux29~4_combout  & (((\reg_file[28][2]~q ) # (!\prif.imemload_id [24])))) # (!\Mux29~4_combout  & (\reg_file[24][2]~q  & ((\prif.imemload_id [24]))))

	.dataa(\Mux29~4_combout ),
	.datab(\reg_file[24][2]~q ),
	.datac(\reg_file[28][2]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux29~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~5 .lut_mask = 16'hE4AA;
defparam \Mux29~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N20
cycloneive_lcell_comb \Mux29~2 (
// Equation(s):
// \Mux29~2_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[22][2]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & ((\reg_file[18][2]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[22][2]~q ),
	.datad(\reg_file[18][2]~q ),
	.cin(gnd),
	.combout(\Mux29~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~2 .lut_mask = 16'hB9A8;
defparam \Mux29~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N15
dffeas \reg_file[30][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][2] .is_wysiwyg = "true";
defparam \reg_file[30][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N14
cycloneive_lcell_comb \Mux29~3 (
// Equation(s):
// \Mux29~3_combout  = (\prif.imemload_id [24] & ((\Mux29~2_combout  & (\reg_file[30][2]~q )) # (!\Mux29~2_combout  & ((\reg_file[26][2]~q ))))) # (!\prif.imemload_id [24] & (\Mux29~2_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux29~2_combout ),
	.datac(\reg_file[30][2]~q ),
	.datad(\reg_file[26][2]~q ),
	.cin(gnd),
	.combout(\Mux29~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~3 .lut_mask = 16'hE6C4;
defparam \Mux29~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N20
cycloneive_lcell_comb \Mux29~6 (
// Equation(s):
// \Mux29~6_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\Mux29~3_combout ))) # (!\prif.imemload_id [22] & (\Mux29~5_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\Mux29~5_combout ),
	.datac(prifimemload_id_22),
	.datad(\Mux29~3_combout ),
	.cin(gnd),
	.combout(\Mux29~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~6 .lut_mask = 16'hF4A4;
defparam \Mux29~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N24
cycloneive_lcell_comb \Mux29~17 (
// Equation(s):
// \Mux29~17_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[13][2]~q ))) # (!\prif.imemload_id [21] & (\reg_file[12][2]~q ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[12][2]~q ),
	.datac(\reg_file[13][2]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux29~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~17 .lut_mask = 16'hFA44;
defparam \Mux29~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N12
cycloneive_lcell_comb \Mux29~18 (
// Equation(s):
// \Mux29~18_combout  = (\prif.imemload_id [22] & ((\Mux29~17_combout  & (\reg_file[15][2]~q )) # (!\Mux29~17_combout  & ((\reg_file[14][2]~q ))))) # (!\prif.imemload_id [22] & (((\Mux29~17_combout ))))

	.dataa(\reg_file[15][2]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[14][2]~q ),
	.datad(\Mux29~17_combout ),
	.cin(gnd),
	.combout(\Mux29~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~18 .lut_mask = 16'hBBC0;
defparam \Mux29~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N15
dffeas \reg_file[6][2] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][2]~67_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][2]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][2] .is_wysiwyg = "true";
defparam \reg_file[6][2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N12
cycloneive_lcell_comb \Mux29~10 (
// Equation(s):
// \Mux29~10_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[5][2]~q )) # (!\prif.imemload_id [21] & ((\reg_file[4][2]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[5][2]~q ),
	.datad(\reg_file[4][2]~q ),
	.cin(gnd),
	.combout(\Mux29~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~10 .lut_mask = 16'hD9C8;
defparam \Mux29~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N14
cycloneive_lcell_comb \Mux29~11 (
// Equation(s):
// \Mux29~11_combout  = (\prif.imemload_id [22] & ((\Mux29~10_combout  & (\reg_file[7][2]~q )) # (!\Mux29~10_combout  & ((\reg_file[6][2]~q ))))) # (!\prif.imemload_id [22] & (((\Mux29~10_combout ))))

	.dataa(\reg_file[7][2]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[6][2]~q ),
	.datad(\Mux29~10_combout ),
	.cin(gnd),
	.combout(\Mux29~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~11 .lut_mask = 16'hBBC0;
defparam \Mux29~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N0
cycloneive_lcell_comb \Mux29~15 (
// Equation(s):
// \Mux29~15_combout  = (\Mux29~14_combout ) # ((\prif.imemload_id [22] & (!\prif.imemload_id [21] & \reg_file[2][2]~q )))

	.dataa(\Mux29~14_combout ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\reg_file[2][2]~q ),
	.cin(gnd),
	.combout(\Mux29~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~15 .lut_mask = 16'hAEAA;
defparam \Mux29~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N10
cycloneive_lcell_comb \Mux29~13 (
// Equation(s):
// \Mux29~13_combout  = (\Mux29~12_combout  & (((\reg_file[11][2]~q ) # (!\prif.imemload_id [21])))) # (!\Mux29~12_combout  & (\reg_file[9][2]~q  & ((\prif.imemload_id [21]))))

	.dataa(\Mux29~12_combout ),
	.datab(\reg_file[9][2]~q ),
	.datac(\reg_file[11][2]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux29~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~13 .lut_mask = 16'hE4AA;
defparam \Mux29~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y25_N18
cycloneive_lcell_comb \Mux29~16 (
// Equation(s):
// \Mux29~16_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\Mux29~13_combout ))) # (!\prif.imemload_id [24] & (\Mux29~15_combout ))))

	.dataa(\Mux29~15_combout ),
	.datab(prifimemload_id_23),
	.datac(\Mux29~13_combout ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux29~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux29~16 .lut_mask = 16'hFC22;
defparam \Mux29~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N30
cycloneive_lcell_comb \Mux27~0 (
// Equation(s):
// \Mux27~0_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][4]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][4]~q )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[25][4]~q ),
	.datad(\reg_file[17][4]~q ),
	.cin(gnd),
	.combout(\Mux27~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~0 .lut_mask = 16'hD9C8;
defparam \Mux27~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y24_N0
cycloneive_lcell_comb \Mux27~1 (
// Equation(s):
// \Mux27~1_combout  = (\prif.imemload_id [23] & ((\Mux27~0_combout  & ((\reg_file[29][4]~q ))) # (!\Mux27~0_combout  & (\reg_file[21][4]~q )))) # (!\prif.imemload_id [23] & (((\Mux27~0_combout ))))

	.dataa(\reg_file[21][4]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[29][4]~q ),
	.datad(\Mux27~0_combout ),
	.cin(gnd),
	.combout(\Mux27~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~1 .lut_mask = 16'hF388;
defparam \Mux27~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N30
cycloneive_lcell_comb \Mux27~7 (
// Equation(s):
// \Mux27~7_combout  = (\prif.imemload_id [24] & ((\reg_file[27][4]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[19][4]~q  & !\prif.imemload_id [23]))))

	.dataa(\reg_file[27][4]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[19][4]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux27~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~7 .lut_mask = 16'hCCB8;
defparam \Mux27~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N14
cycloneive_lcell_comb \Mux27~8 (
// Equation(s):
// \Mux27~8_combout  = (\Mux27~7_combout  & (((\reg_file[31][4]~q ) # (!\prif.imemload_id [23])))) # (!\Mux27~7_combout  & (\reg_file[23][4]~q  & ((\prif.imemload_id [23]))))

	.dataa(\Mux27~7_combout ),
	.datab(\reg_file[23][4]~q ),
	.datac(\reg_file[31][4]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux27~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~8 .lut_mask = 16'hE4AA;
defparam \Mux27~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y34_N23
dffeas \reg_file[16][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][4] .is_wysiwyg = "true";
defparam \reg_file[16][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N22
cycloneive_lcell_comb \Mux27~4 (
// Equation(s):
// \Mux27~4_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[20][4]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[16][4]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][4]~q ),
	.datad(\reg_file[20][4]~q ),
	.cin(gnd),
	.combout(\Mux27~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~4 .lut_mask = 16'hBA98;
defparam \Mux27~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N25
dffeas \reg_file[24][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][4] .is_wysiwyg = "true";
defparam \reg_file[24][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N6
cycloneive_lcell_comb \Mux27~5 (
// Equation(s):
// \Mux27~5_combout  = (\prif.imemload_id [24] & ((\Mux27~4_combout  & (\reg_file[28][4]~q )) # (!\Mux27~4_combout  & ((\reg_file[24][4]~q ))))) # (!\prif.imemload_id [24] & (\Mux27~4_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux27~4_combout ),
	.datac(\reg_file[28][4]~q ),
	.datad(\reg_file[24][4]~q ),
	.cin(gnd),
	.combout(\Mux27~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~5 .lut_mask = 16'hE6C4;
defparam \Mux27~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N28
cycloneive_lcell_comb \Mux27~3 (
// Equation(s):
// \Mux27~3_combout  = (\Mux27~2_combout  & (((\reg_file[30][4]~q )) # (!\prif.imemload_id [24]))) # (!\Mux27~2_combout  & (\prif.imemload_id [24] & (\reg_file[26][4]~q )))

	.dataa(\Mux27~2_combout ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[26][4]~q ),
	.datad(\reg_file[30][4]~q ),
	.cin(gnd),
	.combout(\Mux27~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~3 .lut_mask = 16'hEA62;
defparam \Mux27~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N24
cycloneive_lcell_comb \Mux27~6 (
// Equation(s):
// \Mux27~6_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\Mux27~3_combout ))) # (!\prif.imemload_id [22] & (\Mux27~5_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\Mux27~5_combout ),
	.datac(prifimemload_id_22),
	.datad(\Mux27~3_combout ),
	.cin(gnd),
	.combout(\Mux27~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~6 .lut_mask = 16'hF4A4;
defparam \Mux27~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N20
cycloneive_lcell_comb \reg_file[6][4]~feeder (
// Equation(s):
// \reg_file[6][4]~feeder_combout  = \reg_file_nxt[31][4]~68_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][4]~68_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][4]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][4]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][4]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y27_N21
dffeas \reg_file[6][4] (
	.clk(!CLK),
	.d(\reg_file[6][4]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][4] .is_wysiwyg = "true";
defparam \reg_file[6][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N24
cycloneive_lcell_comb \Mux27~10 (
// Equation(s):
// \Mux27~10_combout  = (\prif.imemload_id [21] & (((\reg_file[5][4]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[4][4]~q  & ((!\prif.imemload_id [22]))))

	.dataa(\reg_file[4][4]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[5][4]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux27~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~10 .lut_mask = 16'hCCE2;
defparam \Mux27~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y25_N24
cycloneive_lcell_comb \Mux27~11 (
// Equation(s):
// \Mux27~11_combout  = (\Mux27~10_combout  & (((\reg_file[7][4]~q ) # (!\prif.imemload_id [22])))) # (!\Mux27~10_combout  & (\reg_file[6][4]~q  & ((\prif.imemload_id [22]))))

	.dataa(\reg_file[6][4]~q ),
	.datab(\Mux27~10_combout ),
	.datac(\reg_file[7][4]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux27~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~11 .lut_mask = 16'hE2CC;
defparam \Mux27~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N20
cycloneive_lcell_comb \Mux27~17 (
// Equation(s):
// \Mux27~17_combout  = (\prif.imemload_id [21] & (((\reg_file[13][4]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[12][4]~q  & ((!\prif.imemload_id [22]))))

	.dataa(\reg_file[12][4]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[13][4]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux27~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~17 .lut_mask = 16'hCCE2;
defparam \Mux27~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N20
cycloneive_lcell_comb \Mux27~18 (
// Equation(s):
// \Mux27~18_combout  = (\prif.imemload_id [22] & ((\Mux27~17_combout  & (\reg_file[15][4]~q )) # (!\Mux27~17_combout  & ((\reg_file[14][4]~q ))))) # (!\prif.imemload_id [22] & (((\Mux27~17_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[15][4]~q ),
	.datac(\reg_file[14][4]~q ),
	.datad(\Mux27~17_combout ),
	.cin(gnd),
	.combout(\Mux27~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~18 .lut_mask = 16'hDDA0;
defparam \Mux27~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y25_N23
dffeas \reg_file[3][4] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][4]~68_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][4]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][4] .is_wysiwyg = "true";
defparam \reg_file[3][4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N22
cycloneive_lcell_comb \Mux27~14 (
// Equation(s):
// \Mux27~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][4]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][4]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][4]~q ),
	.datad(\reg_file[1][4]~q ),
	.cin(gnd),
	.combout(\Mux27~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~14 .lut_mask = 16'hA280;
defparam \Mux27~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N26
cycloneive_lcell_comb \Mux27~15 (
// Equation(s):
// \Mux27~15_combout  = (\Mux27~14_combout ) # ((!\prif.imemload_id [21] & (\prif.imemload_id [22] & \reg_file[2][4]~q )))

	.dataa(prifimemload_id_21),
	.datab(\Mux27~14_combout ),
	.datac(prifimemload_id_22),
	.datad(\reg_file[2][4]~q ),
	.cin(gnd),
	.combout(\Mux27~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~15 .lut_mask = 16'hDCCC;
defparam \Mux27~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N6
cycloneive_lcell_comb \Mux27~13 (
// Equation(s):
// \Mux27~13_combout  = (\Mux27~12_combout  & (((\reg_file[11][4]~q )) # (!\prif.imemload_id [21]))) # (!\Mux27~12_combout  & (\prif.imemload_id [21] & ((\reg_file[9][4]~q ))))

	.dataa(\Mux27~12_combout ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[11][4]~q ),
	.datad(\reg_file[9][4]~q ),
	.cin(gnd),
	.combout(\Mux27~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~13 .lut_mask = 16'hE6A2;
defparam \Mux27~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N28
cycloneive_lcell_comb \Mux27~16 (
// Equation(s):
// \Mux27~16_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\Mux27~13_combout ))) # (!\prif.imemload_id [24] & (\Mux27~15_combout ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux27~15_combout ),
	.datad(\Mux27~13_combout ),
	.cin(gnd),
	.combout(\Mux27~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux27~16 .lut_mask = 16'hDC98;
defparam \Mux27~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N30
cycloneive_lcell_comb \Mux28~7 (
// Equation(s):
// \Mux28~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][3]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][3]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][3]~q ),
	.datad(\reg_file[23][3]~q ),
	.cin(gnd),
	.combout(\Mux28~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~7 .lut_mask = 16'hDC98;
defparam \Mux28~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N26
cycloneive_lcell_comb \Mux28~8 (
// Equation(s):
// \Mux28~8_combout  = (\Mux28~7_combout  & (((\reg_file[31][3]~q )) # (!\prif.imemload_id [24]))) # (!\Mux28~7_combout  & (\prif.imemload_id [24] & ((\reg_file[27][3]~q ))))

	.dataa(\Mux28~7_combout ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[31][3]~q ),
	.datad(\reg_file[27][3]~q ),
	.cin(gnd),
	.combout(\Mux28~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~8 .lut_mask = 16'hE6A2;
defparam \Mux28~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N11
dffeas \reg_file[26][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][3] .is_wysiwyg = "true";
defparam \reg_file[26][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N10
cycloneive_lcell_comb \Mux28~2 (
// Equation(s):
// \Mux28~2_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[26][3]~q ))) # (!\prif.imemload_id [24] & (\reg_file[18][3]~q ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[18][3]~q ),
	.datac(\reg_file[26][3]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux28~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~2 .lut_mask = 16'hFA44;
defparam \Mux28~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N10
cycloneive_lcell_comb \Mux28~3 (
// Equation(s):
// \Mux28~3_combout  = (\prif.imemload_id [23] & ((\Mux28~2_combout  & ((\reg_file[30][3]~q ))) # (!\Mux28~2_combout  & (\reg_file[22][3]~q )))) # (!\prif.imemload_id [23] & (((\Mux28~2_combout ))))

	.dataa(\reg_file[22][3]~q ),
	.datab(prifimemload_id_23),
	.datac(\Mux28~2_combout ),
	.datad(\reg_file[30][3]~q ),
	.cin(gnd),
	.combout(\Mux28~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~3 .lut_mask = 16'hF838;
defparam \Mux28~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N29
dffeas \reg_file[24][3] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][3]~66_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][3]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][3] .is_wysiwyg = "true";
defparam \reg_file[24][3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N28
cycloneive_lcell_comb \Mux28~4 (
// Equation(s):
// \Mux28~4_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[24][3]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & ((\reg_file[16][3]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[24][3]~q ),
	.datad(\reg_file[16][3]~q ),
	.cin(gnd),
	.combout(\Mux28~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~4 .lut_mask = 16'hB9A8;
defparam \Mux28~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N0
cycloneive_lcell_comb \Mux28~5 (
// Equation(s):
// \Mux28~5_combout  = (\prif.imemload_id [23] & ((\Mux28~4_combout  & ((\reg_file[28][3]~q ))) # (!\Mux28~4_combout  & (\reg_file[20][3]~q )))) # (!\prif.imemload_id [23] & (\Mux28~4_combout ))

	.dataa(prifimemload_id_23),
	.datab(\Mux28~4_combout ),
	.datac(\reg_file[20][3]~q ),
	.datad(\reg_file[28][3]~q ),
	.cin(gnd),
	.combout(\Mux28~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~5 .lut_mask = 16'hEC64;
defparam \Mux28~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N8
cycloneive_lcell_comb \Mux28~6 (
// Equation(s):
// \Mux28~6_combout  = (\prif.imemload_id [22] & ((\Mux28~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\Mux28~5_combout  & !\prif.imemload_id [21]))))

	.dataa(\Mux28~3_combout ),
	.datab(\Mux28~5_combout ),
	.datac(prifimemload_id_22),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux28~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~6 .lut_mask = 16'hF0AC;
defparam \Mux28~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N2
cycloneive_lcell_comb \Mux28~0 (
// Equation(s):
// \Mux28~0_combout  = (\prif.imemload_id [23] & (((\reg_file[21][3]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[17][3]~q  & ((!\prif.imemload_id [24]))))

	.dataa(\reg_file[17][3]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[21][3]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux28~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~0 .lut_mask = 16'hCCE2;
defparam \Mux28~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y30_N22
cycloneive_lcell_comb \Mux28~1 (
// Equation(s):
// \Mux28~1_combout  = (\Mux28~0_combout  & (((\reg_file[29][3]~q ) # (!\prif.imemload_id [24])))) # (!\Mux28~0_combout  & (\reg_file[25][3]~q  & ((\prif.imemload_id [24]))))

	.dataa(\reg_file[25][3]~q ),
	.datab(\reg_file[29][3]~q ),
	.datac(\Mux28~0_combout ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux28~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~1 .lut_mask = 16'hCAF0;
defparam \Mux28~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N26
cycloneive_lcell_comb \Mux28~15 (
// Equation(s):
// \Mux28~15_combout  = (\Mux28~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][3]~q  & !\prif.imemload_id [21])))

	.dataa(\Mux28~14_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][3]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux28~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~15 .lut_mask = 16'hAAEA;
defparam \Mux28~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N10
cycloneive_lcell_comb \Mux28~12 (
// Equation(s):
// \Mux28~12_combout  = (\prif.imemload_id [21] & ((\reg_file[5][3]~q ) # ((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (((\reg_file[4][3]~q  & !\prif.imemload_id [22]))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[5][3]~q ),
	.datac(\reg_file[4][3]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux28~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~12 .lut_mask = 16'hAAD8;
defparam \Mux28~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N2
cycloneive_lcell_comb \Mux28~13 (
// Equation(s):
// \Mux28~13_combout  = (\prif.imemload_id [22] & ((\Mux28~12_combout  & ((\reg_file[7][3]~q ))) # (!\Mux28~12_combout  & (\reg_file[6][3]~q )))) # (!\prif.imemload_id [22] & (((\Mux28~12_combout ))))

	.dataa(\reg_file[6][3]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[7][3]~q ),
	.datad(\Mux28~12_combout ),
	.cin(gnd),
	.combout(\Mux28~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~13 .lut_mask = 16'hF388;
defparam \Mux28~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N14
cycloneive_lcell_comb \Mux28~16 (
// Equation(s):
// \Mux28~16_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24]) # (\Mux28~13_combout )))) # (!\prif.imemload_id [23] & (\Mux28~15_combout  & (!\prif.imemload_id [24])))

	.dataa(\Mux28~15_combout ),
	.datab(prifimemload_id_23),
	.datac(prifimemload_id_24),
	.datad(\Mux28~13_combout ),
	.cin(gnd),
	.combout(\Mux28~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~16 .lut_mask = 16'hCEC2;
defparam \Mux28~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N16
cycloneive_lcell_comb \Mux28~10 (
// Equation(s):
// \Mux28~10_combout  = (\prif.imemload_id [22] & (((\reg_file[10][3]~q ) # (\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (\reg_file[8][3]~q  & ((!\prif.imemload_id [21]))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[8][3]~q ),
	.datac(\reg_file[10][3]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux28~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~10 .lut_mask = 16'hAAE4;
defparam \Mux28~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N4
cycloneive_lcell_comb \Mux28~11 (
// Equation(s):
// \Mux28~11_combout  = (\prif.imemload_id [21] & ((\Mux28~10_combout  & (\reg_file[11][3]~q )) # (!\Mux28~10_combout  & ((\reg_file[9][3]~q ))))) # (!\prif.imemload_id [21] & (((\Mux28~10_combout ))))

	.dataa(\reg_file[11][3]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[9][3]~q ),
	.datad(\Mux28~10_combout ),
	.cin(gnd),
	.combout(\Mux28~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~11 .lut_mask = 16'hBBC0;
defparam \Mux28~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N18
cycloneive_lcell_comb \Mux28~17 (
// Equation(s):
// \Mux28~17_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[13][3]~q ))) # (!\prif.imemload_id [21] & (\reg_file[12][3]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[12][3]~q ),
	.datad(\reg_file[13][3]~q ),
	.cin(gnd),
	.combout(\Mux28~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~17 .lut_mask = 16'hDC98;
defparam \Mux28~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N2
cycloneive_lcell_comb \Mux28~18 (
// Equation(s):
// \Mux28~18_combout  = (\Mux28~17_combout  & ((\reg_file[15][3]~q ) # ((!\prif.imemload_id [22])))) # (!\Mux28~17_combout  & (((\reg_file[14][3]~q  & \prif.imemload_id [22]))))

	.dataa(\Mux28~17_combout ),
	.datab(\reg_file[15][3]~q ),
	.datac(\reg_file[14][3]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux28~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux28~18 .lut_mask = 16'hD8AA;
defparam \Mux28~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N18
cycloneive_lcell_comb \Mux23~7 (
// Equation(s):
// \Mux23~7_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[27][8]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[19][8]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][8]~q ),
	.datad(\reg_file[27][8]~q ),
	.cin(gnd),
	.combout(\Mux23~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~7 .lut_mask = 16'hBA98;
defparam \Mux23~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N10
cycloneive_lcell_comb \Mux23~8 (
// Equation(s):
// \Mux23~8_combout  = (\prif.imemload_id [23] & ((\Mux23~7_combout  & ((\reg_file[31][8]~q ))) # (!\Mux23~7_combout  & (\reg_file[23][8]~q )))) # (!\prif.imemload_id [23] & (((\Mux23~7_combout ))))

	.dataa(\reg_file[23][8]~q ),
	.datab(\reg_file[31][8]~q ),
	.datac(prifimemload_id_23),
	.datad(\Mux23~7_combout ),
	.cin(gnd),
	.combout(\Mux23~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~8 .lut_mask = 16'hCFA0;
defparam \Mux23~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N28
cycloneive_lcell_comb \Mux23~2 (
// Equation(s):
// \Mux23~2_combout  = (\prif.imemload_id [23] & ((\reg_file[22][8]~q ) # ((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (((\reg_file[18][8]~q  & !\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[22][8]~q ),
	.datac(\reg_file[18][8]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux23~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~2 .lut_mask = 16'hAAD8;
defparam \Mux23~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N31
dffeas \reg_file[30][8] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][8]~92_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][8] .is_wysiwyg = "true";
defparam \reg_file[30][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N30
cycloneive_lcell_comb \Mux23~3 (
// Equation(s):
// \Mux23~3_combout  = (\prif.imemload_id [24] & ((\Mux23~2_combout  & (\reg_file[30][8]~q )) # (!\Mux23~2_combout  & ((\reg_file[26][8]~q ))))) # (!\prif.imemload_id [24] & (\Mux23~2_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux23~2_combout ),
	.datac(\reg_file[30][8]~q ),
	.datad(\reg_file[26][8]~q ),
	.cin(gnd),
	.combout(\Mux23~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~3 .lut_mask = 16'hE6C4;
defparam \Mux23~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N4
cycloneive_lcell_comb \Mux23~4 (
// Equation(s):
// \Mux23~4_combout  = (\prif.imemload_id [23] & (((\reg_file[20][8]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[16][8]~q  & ((!\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[16][8]~q ),
	.datac(\reg_file[20][8]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux23~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~4 .lut_mask = 16'hAAE4;
defparam \Mux23~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N30
cycloneive_lcell_comb \Mux23~5 (
// Equation(s):
// \Mux23~5_combout  = (\prif.imemload_id [24] & ((\Mux23~4_combout  & ((\reg_file[28][8]~q ))) # (!\Mux23~4_combout  & (\reg_file[24][8]~q )))) # (!\prif.imemload_id [24] & (((\Mux23~4_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[24][8]~q ),
	.datac(\reg_file[28][8]~q ),
	.datad(\Mux23~4_combout ),
	.cin(gnd),
	.combout(\Mux23~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~5 .lut_mask = 16'hF588;
defparam \Mux23~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N8
cycloneive_lcell_comb \Mux23~6 (
// Equation(s):
// \Mux23~6_combout  = (\prif.imemload_id [22] & ((\prif.imemload_id [21]) # ((\Mux23~3_combout )))) # (!\prif.imemload_id [22] & (!\prif.imemload_id [21] & ((\Mux23~5_combout ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\Mux23~3_combout ),
	.datad(\Mux23~5_combout ),
	.cin(gnd),
	.combout(\Mux23~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~6 .lut_mask = 16'hB9A8;
defparam \Mux23~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y28_N22
cycloneive_lcell_comb \reg_file[21][8]~feeder (
// Equation(s):
// \reg_file[21][8]~feeder_combout  = \reg_file_nxt[31][8]~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][8]~92_combout ),
	.cin(gnd),
	.combout(\reg_file[21][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][8]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[21][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y28_N23
dffeas \reg_file[21][8] (
	.clk(!CLK),
	.d(\reg_file[21][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][8] .is_wysiwyg = "true";
defparam \reg_file[21][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N14
cycloneive_lcell_comb \Mux23~0 (
// Equation(s):
// \Mux23~0_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][8]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][8]~q )))))

	.dataa(\reg_file[25][8]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[17][8]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux23~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~0 .lut_mask = 16'hEE30;
defparam \Mux23~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N10
cycloneive_lcell_comb \Mux23~1 (
// Equation(s):
// \Mux23~1_combout  = (\prif.imemload_id [23] & ((\Mux23~0_combout  & ((\reg_file[29][8]~q ))) # (!\Mux23~0_combout  & (\reg_file[21][8]~q )))) # (!\prif.imemload_id [23] & (((\Mux23~0_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[21][8]~q ),
	.datac(\reg_file[29][8]~q ),
	.datad(\Mux23~0_combout ),
	.cin(gnd),
	.combout(\Mux23~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~1 .lut_mask = 16'hF588;
defparam \Mux23~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N8
cycloneive_lcell_comb \Mux23~10 (
// Equation(s):
// \Mux23~10_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[5][8]~q )) # (!\prif.imemload_id [21] & ((\reg_file[4][8]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[5][8]~q ),
	.datad(\reg_file[4][8]~q ),
	.cin(gnd),
	.combout(\Mux23~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~10 .lut_mask = 16'hD9C8;
defparam \Mux23~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N12
cycloneive_lcell_comb \reg_file[7][8]~feeder (
// Equation(s):
// \reg_file[7][8]~feeder_combout  = \reg_file_nxt[31][8]~92_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][8]~92_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[7][8]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[7][8]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[7][8]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y26_N13
dffeas \reg_file[7][8] (
	.clk(!CLK),
	.d(\reg_file[7][8]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][8]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][8] .is_wysiwyg = "true";
defparam \reg_file[7][8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N22
cycloneive_lcell_comb \Mux23~11 (
// Equation(s):
// \Mux23~11_combout  = (\prif.imemload_id [22] & ((\Mux23~10_combout  & ((\reg_file[7][8]~q ))) # (!\Mux23~10_combout  & (\reg_file[6][8]~q )))) # (!\prif.imemload_id [22] & (\Mux23~10_combout ))

	.dataa(prifimemload_id_22),
	.datab(\Mux23~10_combout ),
	.datac(\reg_file[6][8]~q ),
	.datad(\reg_file[7][8]~q ),
	.cin(gnd),
	.combout(\Mux23~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~11 .lut_mask = 16'hEC64;
defparam \Mux23~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N4
cycloneive_lcell_comb \Mux23~17 (
// Equation(s):
// \Mux23~17_combout  = (\prif.imemload_id [21] & (((\reg_file[13][8]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[12][8]~q  & ((!\prif.imemload_id [22]))))

	.dataa(\reg_file[12][8]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[13][8]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux23~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~17 .lut_mask = 16'hCCE2;
defparam \Mux23~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y27_N4
cycloneive_lcell_comb \Mux23~18 (
// Equation(s):
// \Mux23~18_combout  = (\Mux23~17_combout  & (((\reg_file[15][8]~q ) # (!\prif.imemload_id [22])))) # (!\Mux23~17_combout  & (\reg_file[14][8]~q  & (\prif.imemload_id [22])))

	.dataa(\Mux23~17_combout ),
	.datab(\reg_file[14][8]~q ),
	.datac(prifimemload_id_22),
	.datad(\reg_file[15][8]~q ),
	.cin(gnd),
	.combout(\Mux23~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~18 .lut_mask = 16'hEA4A;
defparam \Mux23~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N10
cycloneive_lcell_comb \Mux23~15 (
// Equation(s):
// \Mux23~15_combout  = (\Mux23~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][8]~q  & !\prif.imemload_id [21])))

	.dataa(\Mux23~14_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][8]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux23~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~15 .lut_mask = 16'hAAEA;
defparam \Mux23~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N24
cycloneive_lcell_comb \Mux23~12 (
// Equation(s):
// \Mux23~12_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[10][8]~q ))) # (!\prif.imemload_id [22] & (\reg_file[8][8]~q ))))

	.dataa(\reg_file[8][8]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[10][8]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux23~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~12 .lut_mask = 16'hFC22;
defparam \Mux23~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N14
cycloneive_lcell_comb \Mux23~13 (
// Equation(s):
// \Mux23~13_combout  = (\prif.imemload_id [21] & ((\Mux23~12_combout  & ((\reg_file[11][8]~q ))) # (!\Mux23~12_combout  & (\reg_file[9][8]~q )))) # (!\prif.imemload_id [21] & (((\Mux23~12_combout ))))

	.dataa(\reg_file[9][8]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[11][8]~q ),
	.datad(\Mux23~12_combout ),
	.cin(gnd),
	.combout(\Mux23~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~13 .lut_mask = 16'hF388;
defparam \Mux23~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y26_N28
cycloneive_lcell_comb \Mux23~16 (
// Equation(s):
// \Mux23~16_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\Mux23~13_combout ))) # (!\prif.imemload_id [24] & (\Mux23~15_combout ))))

	.dataa(\Mux23~15_combout ),
	.datab(prifimemload_id_23),
	.datac(prifimemload_id_24),
	.datad(\Mux23~13_combout ),
	.cin(gnd),
	.combout(\Mux23~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux23~16 .lut_mask = 16'hF2C2;
defparam \Mux23~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N12
cycloneive_lcell_comb \Mux24~7 (
// Equation(s):
// \Mux24~7_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\reg_file[23][7]~q )) # (!\prif.imemload_id [23] & ((\reg_file[19][7]~q )))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[23][7]~q ),
	.datac(\reg_file[19][7]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux24~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~7 .lut_mask = 16'hEE50;
defparam \Mux24~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N6
cycloneive_lcell_comb \Mux24~8 (
// Equation(s):
// \Mux24~8_combout  = (\prif.imemload_id [24] & ((\Mux24~7_combout  & ((\reg_file[31][7]~q ))) # (!\Mux24~7_combout  & (\reg_file[27][7]~q )))) # (!\prif.imemload_id [24] & (((\Mux24~7_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[27][7]~q ),
	.datac(\reg_file[31][7]~q ),
	.datad(\Mux24~7_combout ),
	.cin(gnd),
	.combout(\Mux24~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~8 .lut_mask = 16'hF588;
defparam \Mux24~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N22
cycloneive_lcell_comb \reg_file[16][7]~feeder (
// Equation(s):
// \reg_file[16][7]~feeder_combout  = \reg_file_nxt[31][7]~93_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][7]~93_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[16][7]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[16][7]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[16][7]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y30_N23
dffeas \reg_file[16][7] (
	.clk(!CLK),
	.d(\reg_file[16][7]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][7] .is_wysiwyg = "true";
defparam \reg_file[16][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N28
cycloneive_lcell_comb \Mux24~4 (
// Equation(s):
// \Mux24~4_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[24][7]~q )) # (!\prif.imemload_id [24] & ((\reg_file[16][7]~q )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[24][7]~q ),
	.datad(\reg_file[16][7]~q ),
	.cin(gnd),
	.combout(\Mux24~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~4 .lut_mask = 16'hD9C8;
defparam \Mux24~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N18
cycloneive_lcell_comb \Mux24~5 (
// Equation(s):
// \Mux24~5_combout  = (\Mux24~4_combout  & (((\reg_file[28][7]~q ) # (!\prif.imemload_id [23])))) # (!\Mux24~4_combout  & (\reg_file[20][7]~q  & ((\prif.imemload_id [23]))))

	.dataa(\reg_file[20][7]~q ),
	.datab(\Mux24~4_combout ),
	.datac(\reg_file[28][7]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux24~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~5 .lut_mask = 16'hE2CC;
defparam \Mux24~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y30_N1
dffeas \reg_file[18][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][7] .is_wysiwyg = "true";
defparam \reg_file[18][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N0
cycloneive_lcell_comb \Mux24~2 (
// Equation(s):
// \Mux24~2_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[26][7]~q )) # (!\prif.imemload_id [24] & ((\reg_file[18][7]~q )))))

	.dataa(\reg_file[26][7]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[18][7]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux24~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~2 .lut_mask = 16'hEE30;
defparam \Mux24~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N10
cycloneive_lcell_comb \Mux24~3 (
// Equation(s):
// \Mux24~3_combout  = (\prif.imemload_id [23] & ((\Mux24~2_combout  & (\reg_file[30][7]~q )) # (!\Mux24~2_combout  & ((\reg_file[22][7]~q ))))) # (!\prif.imemload_id [23] & (((\Mux24~2_combout ))))

	.dataa(\reg_file[30][7]~q ),
	.datab(prifimemload_id_23),
	.datac(\Mux24~2_combout ),
	.datad(\reg_file[22][7]~q ),
	.cin(gnd),
	.combout(\Mux24~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~3 .lut_mask = 16'hBCB0;
defparam \Mux24~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N8
cycloneive_lcell_comb \Mux24~6 (
// Equation(s):
// \Mux24~6_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\Mux24~3_combout ))) # (!\prif.imemload_id [22] & (\Mux24~5_combout ))))

	.dataa(\Mux24~5_combout ),
	.datab(prifimemload_id_21),
	.datac(\Mux24~3_combout ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux24~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~6 .lut_mask = 16'hFC22;
defparam \Mux24~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N10
cycloneive_lcell_comb \Mux24~0 (
// Equation(s):
// \Mux24~0_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[21][7]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[17][7]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[17][7]~q ),
	.datad(\reg_file[21][7]~q ),
	.cin(gnd),
	.combout(\Mux24~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~0 .lut_mask = 16'hBA98;
defparam \Mux24~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N2
cycloneive_lcell_comb \Mux24~1 (
// Equation(s):
// \Mux24~1_combout  = (\prif.imemload_id [24] & ((\Mux24~0_combout  & ((\reg_file[29][7]~q ))) # (!\Mux24~0_combout  & (\reg_file[25][7]~q )))) # (!\prif.imemload_id [24] & (((\Mux24~0_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[25][7]~q ),
	.datac(\Mux24~0_combout ),
	.datad(\reg_file[29][7]~q ),
	.cin(gnd),
	.combout(\Mux24~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~1 .lut_mask = 16'hF858;
defparam \Mux24~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N28
cycloneive_lcell_comb \Mux24~17 (
// Equation(s):
// \Mux24~17_combout  = (\prif.imemload_id [21] & (((\reg_file[13][7]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[12][7]~q  & ((!\prif.imemload_id [22]))))

	.dataa(\reg_file[12][7]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[13][7]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux24~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~17 .lut_mask = 16'hCCE2;
defparam \Mux24~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N4
cycloneive_lcell_comb \Mux24~18 (
// Equation(s):
// \Mux24~18_combout  = (\prif.imemload_id [22] & ((\Mux24~17_combout  & ((\reg_file[15][7]~q ))) # (!\Mux24~17_combout  & (\reg_file[14][7]~q )))) # (!\prif.imemload_id [22] & (((\Mux24~17_combout ))))

	.dataa(\reg_file[14][7]~q ),
	.datab(\reg_file[15][7]~q ),
	.datac(prifimemload_id_22),
	.datad(\Mux24~17_combout ),
	.cin(gnd),
	.combout(\Mux24~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~18 .lut_mask = 16'hCFA0;
defparam \Mux24~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N0
cycloneive_lcell_comb \Mux24~10 (
// Equation(s):
// \Mux24~10_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[10][7]~q )) # (!\prif.imemload_id [22] & ((\reg_file[8][7]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[10][7]~q ),
	.datad(\reg_file[8][7]~q ),
	.cin(gnd),
	.combout(\Mux24~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~10 .lut_mask = 16'hD9C8;
defparam \Mux24~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N7
dffeas \reg_file[9][7] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][7]~93_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][7]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][7] .is_wysiwyg = "true";
defparam \reg_file[9][7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N6
cycloneive_lcell_comb \Mux24~11 (
// Equation(s):
// \Mux24~11_combout  = (\Mux24~10_combout  & (((\reg_file[11][7]~q )) # (!\prif.imemload_id [21]))) # (!\Mux24~10_combout  & (\prif.imemload_id [21] & (\reg_file[9][7]~q )))

	.dataa(\Mux24~10_combout ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[9][7]~q ),
	.datad(\reg_file[11][7]~q ),
	.cin(gnd),
	.combout(\Mux24~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~11 .lut_mask = 16'hEA62;
defparam \Mux24~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N14
cycloneive_lcell_comb \Mux24~12 (
// Equation(s):
// \Mux24~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][7]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[4][7]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[4][7]~q ),
	.datad(\reg_file[5][7]~q ),
	.cin(gnd),
	.combout(\Mux24~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~12 .lut_mask = 16'hBA98;
defparam \Mux24~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N10
cycloneive_lcell_comb \Mux24~13 (
// Equation(s):
// \Mux24~13_combout  = (\prif.imemload_id [22] & ((\Mux24~12_combout  & ((\reg_file[7][7]~q ))) # (!\Mux24~12_combout  & (\reg_file[6][7]~q )))) # (!\prif.imemload_id [22] & (((\Mux24~12_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[6][7]~q ),
	.datac(\reg_file[7][7]~q ),
	.datad(\Mux24~12_combout ),
	.cin(gnd),
	.combout(\Mux24~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~13 .lut_mask = 16'hF588;
defparam \Mux24~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y33_N10
cycloneive_lcell_comb \Mux24~14 (
// Equation(s):
// \Mux24~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][7]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][7]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][7]~q ),
	.datad(\reg_file[1][7]~q ),
	.cin(gnd),
	.combout(\Mux24~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~14 .lut_mask = 16'hA280;
defparam \Mux24~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N20
cycloneive_lcell_comb \Mux24~15 (
// Equation(s):
// \Mux24~15_combout  = (\Mux24~14_combout ) # ((\reg_file[2][7]~q  & (\prif.imemload_id [22] & !\prif.imemload_id [21])))

	.dataa(\reg_file[2][7]~q ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux24~14_combout ),
	.cin(gnd),
	.combout(\Mux24~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~15 .lut_mask = 16'hFF08;
defparam \Mux24~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N6
cycloneive_lcell_comb \Mux24~16 (
// Equation(s):
// \Mux24~16_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\Mux24~13_combout )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & ((\Mux24~15_combout ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux24~13_combout ),
	.datad(\Mux24~15_combout ),
	.cin(gnd),
	.combout(\Mux24~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux24~16 .lut_mask = 16'hB9A8;
defparam \Mux24~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N24
cycloneive_lcell_comb \Mux25~7 (
// Equation(s):
// \Mux25~7_combout  = (\prif.imemload_id [24] & ((\reg_file[27][6]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[19][6]~q  & !\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[27][6]~q ),
	.datac(\reg_file[19][6]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux25~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~7 .lut_mask = 16'hAAD8;
defparam \Mux25~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N18
cycloneive_lcell_comb \Mux25~8 (
// Equation(s):
// \Mux25~8_combout  = (\Mux25~7_combout  & ((\reg_file[31][6]~q ) # ((!\prif.imemload_id [23])))) # (!\Mux25~7_combout  & (((\reg_file[23][6]~q  & \prif.imemload_id [23]))))

	.dataa(\Mux25~7_combout ),
	.datab(\reg_file[31][6]~q ),
	.datac(\reg_file[23][6]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux25~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~8 .lut_mask = 16'hD8AA;
defparam \Mux25~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y32_N11
dffeas \reg_file[20][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][6] .is_wysiwyg = "true";
defparam \reg_file[20][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N10
cycloneive_lcell_comb \Mux25~4 (
// Equation(s):
// \Mux25~4_combout  = (\prif.imemload_id [23] & (((\reg_file[20][6]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[16][6]~q  & ((!\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[16][6]~q ),
	.datac(\reg_file[20][6]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux25~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~4 .lut_mask = 16'hAAE4;
defparam \Mux25~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N28
cycloneive_lcell_comb \Mux25~5 (
// Equation(s):
// \Mux25~5_combout  = (\prif.imemload_id [24] & ((\Mux25~4_combout  & ((\reg_file[28][6]~q ))) # (!\Mux25~4_combout  & (\reg_file[24][6]~q )))) # (!\prif.imemload_id [24] & (((\Mux25~4_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[24][6]~q ),
	.datac(\reg_file[28][6]~q ),
	.datad(\Mux25~4_combout ),
	.cin(gnd),
	.combout(\Mux25~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~5 .lut_mask = 16'hF588;
defparam \Mux25~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y30_N13
dffeas \reg_file[30][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][6] .is_wysiwyg = "true";
defparam \reg_file[30][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N12
cycloneive_lcell_comb \Mux25~3 (
// Equation(s):
// \Mux25~3_combout  = (\Mux25~2_combout  & (((\reg_file[30][6]~q ) # (!\prif.imemload_id [24])))) # (!\Mux25~2_combout  & (\reg_file[26][6]~q  & ((\prif.imemload_id [24]))))

	.dataa(\Mux25~2_combout ),
	.datab(\reg_file[26][6]~q ),
	.datac(\reg_file[30][6]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux25~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~3 .lut_mask = 16'hE4AA;
defparam \Mux25~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N4
cycloneive_lcell_comb \Mux25~6 (
// Equation(s):
// \Mux25~6_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21]) # (\Mux25~3_combout )))) # (!\prif.imemload_id [22] & (\Mux25~5_combout  & (!\prif.imemload_id [21])))

	.dataa(\Mux25~5_combout ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux25~3_combout ),
	.cin(gnd),
	.combout(\Mux25~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~6 .lut_mask = 16'hCEC2;
defparam \Mux25~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y29_N19
dffeas \reg_file[21][6] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][6]~80_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][6]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][6] .is_wysiwyg = "true";
defparam \reg_file[21][6] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N4
cycloneive_lcell_comb \Mux25~0 (
// Equation(s):
// \Mux25~0_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][6]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][6]~q )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[25][6]~q ),
	.datad(\reg_file[17][6]~q ),
	.cin(gnd),
	.combout(\Mux25~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~0 .lut_mask = 16'hD9C8;
defparam \Mux25~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N18
cycloneive_lcell_comb \Mux25~1 (
// Equation(s):
// \Mux25~1_combout  = (\prif.imemload_id [23] & ((\Mux25~0_combout  & (\reg_file[29][6]~q )) # (!\Mux25~0_combout  & ((\reg_file[21][6]~q ))))) # (!\prif.imemload_id [23] & (((\Mux25~0_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[29][6]~q ),
	.datac(\reg_file[21][6]~q ),
	.datad(\Mux25~0_combout ),
	.cin(gnd),
	.combout(\Mux25~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~1 .lut_mask = 16'hDDA0;
defparam \Mux25~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N2
cycloneive_lcell_comb \Mux25~17 (
// Equation(s):
// \Mux25~17_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[13][6]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[12][6]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[12][6]~q ),
	.datad(\reg_file[13][6]~q ),
	.cin(gnd),
	.combout(\Mux25~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~17 .lut_mask = 16'hBA98;
defparam \Mux25~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N6
cycloneive_lcell_comb \Mux25~18 (
// Equation(s):
// \Mux25~18_combout  = (\prif.imemload_id [22] & ((\Mux25~17_combout  & (\reg_file[15][6]~q )) # (!\Mux25~17_combout  & ((\reg_file[14][6]~q ))))) # (!\prif.imemload_id [22] & (((\Mux25~17_combout ))))

	.dataa(\reg_file[15][6]~q ),
	.datab(\reg_file[14][6]~q ),
	.datac(prifimemload_id_22),
	.datad(\Mux25~17_combout ),
	.cin(gnd),
	.combout(\Mux25~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~18 .lut_mask = 16'hAFC0;
defparam \Mux25~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N8
cycloneive_lcell_comb \Mux25~12 (
// Equation(s):
// \Mux25~12_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[10][6]~q )) # (!\prif.imemload_id [22] & ((\reg_file[8][6]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[10][6]~q ),
	.datad(\reg_file[8][6]~q ),
	.cin(gnd),
	.combout(\Mux25~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~12 .lut_mask = 16'hD9C8;
defparam \Mux25~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N8
cycloneive_lcell_comb \Mux25~13 (
// Equation(s):
// \Mux25~13_combout  = (\prif.imemload_id [21] & ((\Mux25~12_combout  & (\reg_file[11][6]~q )) # (!\Mux25~12_combout  & ((\reg_file[9][6]~q ))))) # (!\prif.imemload_id [21] & (((\Mux25~12_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[11][6]~q ),
	.datac(\reg_file[9][6]~q ),
	.datad(\Mux25~12_combout ),
	.cin(gnd),
	.combout(\Mux25~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~13 .lut_mask = 16'hDDA0;
defparam \Mux25~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N22
cycloneive_lcell_comb \Mux25~14 (
// Equation(s):
// \Mux25~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][6]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][6]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[1][6]~q ),
	.datad(\reg_file[3][6]~q ),
	.cin(gnd),
	.combout(\Mux25~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~14 .lut_mask = 16'hA820;
defparam \Mux25~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N20
cycloneive_lcell_comb \Mux25~15 (
// Equation(s):
// \Mux25~15_combout  = (\Mux25~14_combout ) # ((!\prif.imemload_id [21] & (\prif.imemload_id [22] & \reg_file[2][6]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][6]~q ),
	.datad(\Mux25~14_combout ),
	.cin(gnd),
	.combout(\Mux25~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~15 .lut_mask = 16'hFF40;
defparam \Mux25~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N10
cycloneive_lcell_comb \Mux25~16 (
// Equation(s):
// \Mux25~16_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\Mux25~13_combout )) # (!\prif.imemload_id [24] & ((\Mux25~15_combout )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux25~13_combout ),
	.datad(\Mux25~15_combout ),
	.cin(gnd),
	.combout(\Mux25~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~16 .lut_mask = 16'hD9C8;
defparam \Mux25~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N6
cycloneive_lcell_comb \Mux25~10 (
// Equation(s):
// \Mux25~10_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[5][6]~q ))) # (!\prif.imemload_id [21] & (\reg_file[4][6]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[4][6]~q ),
	.datad(\reg_file[5][6]~q ),
	.cin(gnd),
	.combout(\Mux25~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~10 .lut_mask = 16'hDC98;
defparam \Mux25~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N16
cycloneive_lcell_comb \Mux25~11 (
// Equation(s):
// \Mux25~11_combout  = (\Mux25~10_combout  & ((\reg_file[7][6]~q ) # ((!\prif.imemload_id [22])))) # (!\Mux25~10_combout  & (((\reg_file[6][6]~q  & \prif.imemload_id [22]))))

	.dataa(\reg_file[7][6]~q ),
	.datab(\Mux25~10_combout ),
	.datac(\reg_file[6][6]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux25~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux25~11 .lut_mask = 16'hB8CC;
defparam \Mux25~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N4
cycloneive_lcell_comb \Mux26~0 (
// Equation(s):
// \Mux26~0_combout  = (\prif.imemload_id [23] & ((\reg_file[21][5]~q ) # ((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (((\reg_file[17][5]~q  & !\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[21][5]~q ),
	.datac(\reg_file[17][5]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux26~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~0 .lut_mask = 16'hAAD8;
defparam \Mux26~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N30
cycloneive_lcell_comb \Mux26~1 (
// Equation(s):
// \Mux26~1_combout  = (\prif.imemload_id [24] & ((\Mux26~0_combout  & (\reg_file[29][5]~q )) # (!\Mux26~0_combout  & ((\reg_file[25][5]~q ))))) # (!\prif.imemload_id [24] & (((\Mux26~0_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[29][5]~q ),
	.datac(\reg_file[25][5]~q ),
	.datad(\Mux26~0_combout ),
	.cin(gnd),
	.combout(\Mux26~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~1 .lut_mask = 16'hDDA0;
defparam \Mux26~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N2
cycloneive_lcell_comb \Mux26~7 (
// Equation(s):
// \Mux26~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][5]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][5]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][5]~q ),
	.datad(\reg_file[23][5]~q ),
	.cin(gnd),
	.combout(\Mux26~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~7 .lut_mask = 16'hDC98;
defparam \Mux26~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N2
cycloneive_lcell_comb \Mux26~8 (
// Equation(s):
// \Mux26~8_combout  = (\prif.imemload_id [24] & ((\Mux26~7_combout  & ((\reg_file[31][5]~q ))) # (!\Mux26~7_combout  & (\reg_file[27][5]~q )))) # (!\prif.imemload_id [24] & (((\Mux26~7_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[27][5]~q ),
	.datac(\reg_file[31][5]~q ),
	.datad(\Mux26~7_combout ),
	.cin(gnd),
	.combout(\Mux26~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~8 .lut_mask = 16'hF588;
defparam \Mux26~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N18
cycloneive_lcell_comb \Mux26~4 (
// Equation(s):
// \Mux26~4_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[24][5]~q ))) # (!\prif.imemload_id [24] & (\reg_file[16][5]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][5]~q ),
	.datad(\reg_file[24][5]~q ),
	.cin(gnd),
	.combout(\Mux26~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~4 .lut_mask = 16'hDC98;
defparam \Mux26~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y34_N27
dffeas \reg_file[28][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][5] .is_wysiwyg = "true";
defparam \reg_file[28][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N26
cycloneive_lcell_comb \Mux26~5 (
// Equation(s):
// \Mux26~5_combout  = (\Mux26~4_combout  & (((\reg_file[28][5]~q ) # (!\prif.imemload_id [23])))) # (!\Mux26~4_combout  & (\reg_file[20][5]~q  & ((\prif.imemload_id [23]))))

	.dataa(\reg_file[20][5]~q ),
	.datab(\Mux26~4_combout ),
	.datac(\reg_file[28][5]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux26~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~5 .lut_mask = 16'hE2CC;
defparam \Mux26~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N24
cycloneive_lcell_comb \reg_file[22][5]~feeder (
// Equation(s):
// \reg_file[22][5]~feeder_combout  = \reg_file_nxt[31][5]~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][5]~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[22][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][5]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[22][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N25
dffeas \reg_file[22][5] (
	.clk(!CLK),
	.d(\reg_file[22][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][5] .is_wysiwyg = "true";
defparam \reg_file[22][5] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N13
dffeas \reg_file[18][5] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][5]~72_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][5] .is_wysiwyg = "true";
defparam \reg_file[18][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N14
cycloneive_lcell_comb \Mux26~2 (
// Equation(s):
// \Mux26~2_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[26][5]~q )) # (!\prif.imemload_id [24] & ((\reg_file[18][5]~q )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[26][5]~q ),
	.datad(\reg_file[18][5]~q ),
	.cin(gnd),
	.combout(\Mux26~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~2 .lut_mask = 16'hD9C8;
defparam \Mux26~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N26
cycloneive_lcell_comb \Mux26~3 (
// Equation(s):
// \Mux26~3_combout  = (\prif.imemload_id [23] & ((\Mux26~2_combout  & ((\reg_file[30][5]~q ))) # (!\Mux26~2_combout  & (\reg_file[22][5]~q )))) # (!\prif.imemload_id [23] & (((\Mux26~2_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[22][5]~q ),
	.datac(\reg_file[30][5]~q ),
	.datad(\Mux26~2_combout ),
	.cin(gnd),
	.combout(\Mux26~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~3 .lut_mask = 16'hF588;
defparam \Mux26~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y28_N4
cycloneive_lcell_comb \Mux26~6 (
// Equation(s):
// \Mux26~6_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\Mux26~3_combout ))) # (!\prif.imemload_id [22] & (\Mux26~5_combout ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux26~5_combout ),
	.datad(\Mux26~3_combout ),
	.cin(gnd),
	.combout(\Mux26~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~6 .lut_mask = 16'hDC98;
defparam \Mux26~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N26
cycloneive_lcell_comb \reg_file[2][5]~feeder (
// Equation(s):
// \reg_file[2][5]~feeder_combout  = \reg_file_nxt[31][5]~72_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][5]~72_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[2][5]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[2][5]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[2][5]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y28_N27
dffeas \reg_file[2][5] (
	.clk(!CLK),
	.d(\reg_file[2][5]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][5]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][5] .is_wysiwyg = "true";
defparam \reg_file[2][5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N2
cycloneive_lcell_comb \Mux26~14 (
// Equation(s):
// \Mux26~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][5]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][5]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[3][5]~q ),
	.datad(\reg_file[1][5]~q ),
	.cin(gnd),
	.combout(\Mux26~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~14 .lut_mask = 16'hC480;
defparam \Mux26~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N28
cycloneive_lcell_comb \Mux26~15 (
// Equation(s):
// \Mux26~15_combout  = (\Mux26~14_combout ) # ((!\prif.imemload_id [21] & (\prif.imemload_id [22] & \reg_file[2][5]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][5]~q ),
	.datad(\Mux26~14_combout ),
	.cin(gnd),
	.combout(\Mux26~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~15 .lut_mask = 16'hFF40;
defparam \Mux26~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N4
cycloneive_lcell_comb \Mux26~12 (
// Equation(s):
// \Mux26~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][5]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[4][5]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[4][5]~q ),
	.datad(\reg_file[5][5]~q ),
	.cin(gnd),
	.combout(\Mux26~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~12 .lut_mask = 16'hBA98;
defparam \Mux26~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N30
cycloneive_lcell_comb \Mux26~13 (
// Equation(s):
// \Mux26~13_combout  = (\Mux26~12_combout  & (((\reg_file[7][5]~q ) # (!\prif.imemload_id [22])))) # (!\Mux26~12_combout  & (\reg_file[6][5]~q  & ((\prif.imemload_id [22]))))

	.dataa(\reg_file[6][5]~q ),
	.datab(\Mux26~12_combout ),
	.datac(\reg_file[7][5]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux26~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~13 .lut_mask = 16'hE2CC;
defparam \Mux26~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N6
cycloneive_lcell_comb \Mux26~16 (
// Equation(s):
// \Mux26~16_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24]) # (\Mux26~13_combout )))) # (!\prif.imemload_id [23] & (\Mux26~15_combout  & (!\prif.imemload_id [24])))

	.dataa(prifimemload_id_23),
	.datab(\Mux26~15_combout ),
	.datac(prifimemload_id_24),
	.datad(\Mux26~13_combout ),
	.cin(gnd),
	.combout(\Mux26~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~16 .lut_mask = 16'hAEA4;
defparam \Mux26~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N8
cycloneive_lcell_comb \Mux26~17 (
// Equation(s):
// \Mux26~17_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[13][5]~q ))) # (!\prif.imemload_id [21] & (\reg_file[12][5]~q ))))

	.dataa(\reg_file[12][5]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[13][5]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux26~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~17 .lut_mask = 16'hFC22;
defparam \Mux26~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y28_N0
cycloneive_lcell_comb \Mux26~18 (
// Equation(s):
// \Mux26~18_combout  = (\Mux26~17_combout  & ((\reg_file[15][5]~q ) # ((!\prif.imemload_id [22])))) # (!\Mux26~17_combout  & (((\reg_file[14][5]~q  & \prif.imemload_id [22]))))

	.dataa(\Mux26~17_combout ),
	.datab(\reg_file[15][5]~q ),
	.datac(\reg_file[14][5]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux26~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~18 .lut_mask = 16'hD8AA;
defparam \Mux26~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N4
cycloneive_lcell_comb \Mux26~10 (
// Equation(s):
// \Mux26~10_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[10][5]~q )) # (!\prif.imemload_id [22] & ((\reg_file[8][5]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[10][5]~q ),
	.datad(\reg_file[8][5]~q ),
	.cin(gnd),
	.combout(\Mux26~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~10 .lut_mask = 16'hD9C8;
defparam \Mux26~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N16
cycloneive_lcell_comb \Mux26~11 (
// Equation(s):
// \Mux26~11_combout  = (\prif.imemload_id [21] & ((\Mux26~10_combout  & ((\reg_file[11][5]~q ))) # (!\Mux26~10_combout  & (\reg_file[9][5]~q )))) # (!\prif.imemload_id [21] & (\Mux26~10_combout ))

	.dataa(prifimemload_id_21),
	.datab(\Mux26~10_combout ),
	.datac(\reg_file[9][5]~q ),
	.datad(\reg_file[11][5]~q ),
	.cin(gnd),
	.combout(\Mux26~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux26~11 .lut_mask = 16'hEC64;
defparam \Mux26~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y26_N31
dffeas \reg_file[19][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][16] .is_wysiwyg = "true";
defparam \reg_file[19][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N30
cycloneive_lcell_comb \Mux15~7 (
// Equation(s):
// \Mux15~7_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[27][16]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[19][16]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][16]~q ),
	.datad(\reg_file[27][16]~q ),
	.cin(gnd),
	.combout(\Mux15~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~7 .lut_mask = 16'hBA98;
defparam \Mux15~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N26
cycloneive_lcell_comb \Mux15~8 (
// Equation(s):
// \Mux15~8_combout  = (\prif.imemload_id [23] & ((\Mux15~7_combout  & (\reg_file[31][16]~q )) # (!\Mux15~7_combout  & ((\reg_file[23][16]~q ))))) # (!\prif.imemload_id [23] & (((\Mux15~7_combout ))))

	.dataa(\reg_file[31][16]~q ),
	.datab(\reg_file[23][16]~q ),
	.datac(prifimemload_id_23),
	.datad(\Mux15~7_combout ),
	.cin(gnd),
	.combout(\Mux15~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~8 .lut_mask = 16'hAFC0;
defparam \Mux15~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N30
cycloneive_lcell_comb \reg_file[21][16]~feeder (
// Equation(s):
// \reg_file[21][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][16]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[21][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[21][16]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[21][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y31_N31
dffeas \reg_file[21][16] (
	.clk(!CLK),
	.d(\reg_file[21][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~15_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[21][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[21][16] .is_wysiwyg = "true";
defparam \reg_file[21][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N22
cycloneive_lcell_comb \Mux15~0 (
// Equation(s):
// \Mux15~0_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[25][16]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & ((\reg_file[17][16]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[25][16]~q ),
	.datad(\reg_file[17][16]~q ),
	.cin(gnd),
	.combout(\Mux15~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~0 .lut_mask = 16'hB9A8;
defparam \Mux15~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N26
cycloneive_lcell_comb \Mux15~1 (
// Equation(s):
// \Mux15~1_combout  = (\prif.imemload_id [23] & ((\Mux15~0_combout  & ((\reg_file[29][16]~q ))) # (!\Mux15~0_combout  & (\reg_file[21][16]~q )))) # (!\prif.imemload_id [23] & (((\Mux15~0_combout ))))

	.dataa(\reg_file[21][16]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[29][16]~q ),
	.datad(\Mux15~0_combout ),
	.cin(gnd),
	.combout(\Mux15~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~1 .lut_mask = 16'hF388;
defparam \Mux15~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N27
dffeas \reg_file[26][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][16] .is_wysiwyg = "true";
defparam \reg_file[26][16] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y30_N17
dffeas \reg_file[18][16] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][16]~85_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][16] .is_wysiwyg = "true";
defparam \reg_file[18][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N16
cycloneive_lcell_comb \Mux15~2 (
// Equation(s):
// \Mux15~2_combout  = (\prif.imemload_id [23] & ((\reg_file[22][16]~q ) # ((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (((\reg_file[18][16]~q  & !\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[22][16]~q ),
	.datac(\reg_file[18][16]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux15~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~2 .lut_mask = 16'hAAD8;
defparam \Mux15~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N30
cycloneive_lcell_comb \Mux15~3 (
// Equation(s):
// \Mux15~3_combout  = (\prif.imemload_id [24] & ((\Mux15~2_combout  & (\reg_file[30][16]~q )) # (!\Mux15~2_combout  & ((\reg_file[26][16]~q ))))) # (!\prif.imemload_id [24] & (((\Mux15~2_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[30][16]~q ),
	.datac(\reg_file[26][16]~q ),
	.datad(\Mux15~2_combout ),
	.cin(gnd),
	.combout(\Mux15~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~3 .lut_mask = 16'hDDA0;
defparam \Mux15~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N20
cycloneive_lcell_comb \Mux15~4 (
// Equation(s):
// \Mux15~4_combout  = (\prif.imemload_id [23] & (((\reg_file[20][16]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[16][16]~q  & ((!\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[16][16]~q ),
	.datac(\reg_file[20][16]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux15~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~4 .lut_mask = 16'hAAE4;
defparam \Mux15~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N18
cycloneive_lcell_comb \Mux15~5 (
// Equation(s):
// \Mux15~5_combout  = (\prif.imemload_id [24] & ((\Mux15~4_combout  & ((\reg_file[28][16]~q ))) # (!\Mux15~4_combout  & (\reg_file[24][16]~q )))) # (!\prif.imemload_id [24] & (((\Mux15~4_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[24][16]~q ),
	.datac(\reg_file[28][16]~q ),
	.datad(\Mux15~4_combout ),
	.cin(gnd),
	.combout(\Mux15~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~5 .lut_mask = 16'hF588;
defparam \Mux15~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N28
cycloneive_lcell_comb \Mux15~6 (
// Equation(s):
// \Mux15~6_combout  = (\prif.imemload_id [22] & ((\Mux15~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((!\prif.imemload_id [21] & \Mux15~5_combout ))))

	.dataa(\Mux15~3_combout ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux15~5_combout ),
	.cin(gnd),
	.combout(\Mux15~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~6 .lut_mask = 16'hCBC8;
defparam \Mux15~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N24
cycloneive_lcell_comb \Mux15~17 (
// Equation(s):
// \Mux15~17_combout  = (\prif.imemload_id [21] & (((\reg_file[13][16]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[12][16]~q  & ((!\prif.imemload_id [22]))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[12][16]~q ),
	.datac(\reg_file[13][16]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux15~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~17 .lut_mask = 16'hAAE4;
defparam \Mux15~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N0
cycloneive_lcell_comb \Mux15~18 (
// Equation(s):
// \Mux15~18_combout  = (\prif.imemload_id [22] & ((\Mux15~17_combout  & ((\reg_file[15][16]~q ))) # (!\Mux15~17_combout  & (\reg_file[14][16]~q )))) # (!\prif.imemload_id [22] & (\Mux15~17_combout ))

	.dataa(prifimemload_id_22),
	.datab(\Mux15~17_combout ),
	.datac(\reg_file[14][16]~q ),
	.datad(\reg_file[15][16]~q ),
	.cin(gnd),
	.combout(\Mux15~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~18 .lut_mask = 16'hEC64;
defparam \Mux15~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N4
cycloneive_lcell_comb \Mux15~13 (
// Equation(s):
// \Mux15~13_combout  = (\Mux15~12_combout  & ((\reg_file[11][16]~q ) # ((!\prif.imemload_id [21])))) # (!\Mux15~12_combout  & (((\prif.imemload_id [21] & \reg_file[9][16]~q ))))

	.dataa(\Mux15~12_combout ),
	.datab(\reg_file[11][16]~q ),
	.datac(prifimemload_id_21),
	.datad(\reg_file[9][16]~q ),
	.cin(gnd),
	.combout(\Mux15~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~13 .lut_mask = 16'hDA8A;
defparam \Mux15~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N22
cycloneive_lcell_comb \reg_file[3][16]~feeder (
// Equation(s):
// \reg_file[3][16]~feeder_combout  = \reg_file_nxt[31][16]~85_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][16]~85_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[3][16]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[3][16]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[3][16]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N23
dffeas \reg_file[3][16] (
	.clk(!CLK),
	.d(\reg_file[3][16]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][16]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][16] .is_wysiwyg = "true";
defparam \reg_file[3][16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N10
cycloneive_lcell_comb \Mux15~14 (
// Equation(s):
// \Mux15~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][16]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][16]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][16]~q ),
	.datad(\reg_file[1][16]~q ),
	.cin(gnd),
	.combout(\Mux15~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~14 .lut_mask = 16'hA280;
defparam \Mux15~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N6
cycloneive_lcell_comb \Mux15~15 (
// Equation(s):
// \Mux15~15_combout  = (\Mux15~14_combout ) # ((\prif.imemload_id [22] & (!\prif.imemload_id [21] & \reg_file[2][16]~q )))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[2][16]~q ),
	.datad(\Mux15~14_combout ),
	.cin(gnd),
	.combout(\Mux15~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~15 .lut_mask = 16'hFF20;
defparam \Mux15~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N26
cycloneive_lcell_comb \Mux15~16 (
// Equation(s):
// \Mux15~16_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\Mux15~13_combout )) # (!\prif.imemload_id [24] & ((\Mux15~15_combout )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux15~13_combout ),
	.datad(\Mux15~15_combout ),
	.cin(gnd),
	.combout(\Mux15~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~16 .lut_mask = 16'hD9C8;
defparam \Mux15~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N28
cycloneive_lcell_comb \Mux15~10 (
// Equation(s):
// \Mux15~10_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[5][16]~q )) # (!\prif.imemload_id [21] & ((\reg_file[4][16]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[5][16]~q ),
	.datad(\reg_file[4][16]~q ),
	.cin(gnd),
	.combout(\Mux15~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~10 .lut_mask = 16'hD9C8;
defparam \Mux15~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N8
cycloneive_lcell_comb \Mux15~11 (
// Equation(s):
// \Mux15~11_combout  = (\Mux15~10_combout  & (((\reg_file[7][16]~q )) # (!\prif.imemload_id [22]))) # (!\Mux15~10_combout  & (\prif.imemload_id [22] & (\reg_file[6][16]~q )))

	.dataa(\Mux15~10_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[6][16]~q ),
	.datad(\reg_file[7][16]~q ),
	.cin(gnd),
	.combout(\Mux15~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux15~11 .lut_mask = 16'hEA62;
defparam \Mux15~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N18
cycloneive_lcell_comb \Mux16~0 (
// Equation(s):
// \Mux16~0_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[21][15]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[17][15]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[17][15]~q ),
	.datad(\reg_file[21][15]~q ),
	.cin(gnd),
	.combout(\Mux16~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~0 .lut_mask = 16'hBA98;
defparam \Mux16~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N16
cycloneive_lcell_comb \Mux16~1 (
// Equation(s):
// \Mux16~1_combout  = (\Mux16~0_combout  & ((\reg_file[29][15]~q ) # ((!\prif.imemload_id [24])))) # (!\Mux16~0_combout  & (((\prif.imemload_id [24] & \reg_file[25][15]~q ))))

	.dataa(\Mux16~0_combout ),
	.datab(\reg_file[29][15]~q ),
	.datac(prifimemload_id_24),
	.datad(\reg_file[25][15]~q ),
	.cin(gnd),
	.combout(\Mux16~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~1 .lut_mask = 16'hDA8A;
defparam \Mux16~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N12
cycloneive_lcell_comb \Mux16~7 (
// Equation(s):
// \Mux16~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][15]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][15]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][15]~q ),
	.datad(\reg_file[23][15]~q ),
	.cin(gnd),
	.combout(\Mux16~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~7 .lut_mask = 16'hDC98;
defparam \Mux16~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N20
cycloneive_lcell_comb \Mux16~8 (
// Equation(s):
// \Mux16~8_combout  = (\prif.imemload_id [24] & ((\Mux16~7_combout  & ((\reg_file[31][15]~q ))) # (!\Mux16~7_combout  & (\reg_file[27][15]~q )))) # (!\prif.imemload_id [24] & (((\Mux16~7_combout ))))

	.dataa(\reg_file[27][15]~q ),
	.datab(\reg_file[31][15]~q ),
	.datac(prifimemload_id_24),
	.datad(\Mux16~7_combout ),
	.cin(gnd),
	.combout(\Mux16~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~8 .lut_mask = 16'hCFA0;
defparam \Mux16~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N2
cycloneive_lcell_comb \Mux16~2 (
// Equation(s):
// \Mux16~2_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[26][15]~q ))) # (!\prif.imemload_id [24] & (\reg_file[18][15]~q ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[18][15]~q ),
	.datac(\reg_file[26][15]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux16~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~2 .lut_mask = 16'hFA44;
defparam \Mux16~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N28
cycloneive_lcell_comb \Mux16~3 (
// Equation(s):
// \Mux16~3_combout  = (\prif.imemload_id [23] & ((\Mux16~2_combout  & (\reg_file[30][15]~q )) # (!\Mux16~2_combout  & ((\reg_file[22][15]~q ))))) # (!\prif.imemload_id [23] & (((\Mux16~2_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[30][15]~q ),
	.datac(\reg_file[22][15]~q ),
	.datad(\Mux16~2_combout ),
	.cin(gnd),
	.combout(\Mux16~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~3 .lut_mask = 16'hDDA0;
defparam \Mux16~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N10
cycloneive_lcell_comb \Mux16~4 (
// Equation(s):
// \Mux16~4_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[24][15]~q ))) # (!\prif.imemload_id [24] & (\reg_file[16][15]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][15]~q ),
	.datad(\reg_file[24][15]~q ),
	.cin(gnd),
	.combout(\Mux16~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~4 .lut_mask = 16'hDC98;
defparam \Mux16~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N4
cycloneive_lcell_comb \Mux16~5 (
// Equation(s):
// \Mux16~5_combout  = (\Mux16~4_combout  & (((\reg_file[28][15]~q ) # (!\prif.imemload_id [23])))) # (!\Mux16~4_combout  & (\reg_file[20][15]~q  & ((\prif.imemload_id [23]))))

	.dataa(\reg_file[20][15]~q ),
	.datab(\Mux16~4_combout ),
	.datac(\reg_file[28][15]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux16~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~5 .lut_mask = 16'hE2CC;
defparam \Mux16~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y24_N0
cycloneive_lcell_comb \Mux16~6 (
// Equation(s):
// \Mux16~6_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\Mux16~3_combout )) # (!\prif.imemload_id [22] & ((\Mux16~5_combout )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux16~3_combout ),
	.datad(\Mux16~5_combout ),
	.cin(gnd),
	.combout(\Mux16~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~6 .lut_mask = 16'hD9C8;
defparam \Mux16~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N12
cycloneive_lcell_comb \Mux16~17 (
// Equation(s):
// \Mux16~17_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[13][15]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & ((\reg_file[12][15]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[13][15]~q ),
	.datad(\reg_file[12][15]~q ),
	.cin(gnd),
	.combout(\Mux16~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~17 .lut_mask = 16'hB9A8;
defparam \Mux16~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N0
cycloneive_lcell_comb \Mux16~18 (
// Equation(s):
// \Mux16~18_combout  = (\Mux16~17_combout  & (((\reg_file[15][15]~q ) # (!\prif.imemload_id [22])))) # (!\Mux16~17_combout  & (\reg_file[14][15]~q  & (\prif.imemload_id [22])))

	.dataa(\Mux16~17_combout ),
	.datab(\reg_file[14][15]~q ),
	.datac(prifimemload_id_22),
	.datad(\reg_file[15][15]~q ),
	.cin(gnd),
	.combout(\Mux16~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~18 .lut_mask = 16'hEA4A;
defparam \Mux16~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N16
cycloneive_lcell_comb \Mux16~10 (
// Equation(s):
// \Mux16~10_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[10][15]~q ))) # (!\prif.imemload_id [22] & (\reg_file[8][15]~q ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[8][15]~q ),
	.datac(\reg_file[10][15]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux16~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~10 .lut_mask = 16'hFA44;
defparam \Mux16~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N14
cycloneive_lcell_comb \Mux16~11 (
// Equation(s):
// \Mux16~11_combout  = (\Mux16~10_combout  & ((\reg_file[11][15]~q ) # ((!\prif.imemload_id [21])))) # (!\Mux16~10_combout  & (((\reg_file[9][15]~q  & \prif.imemload_id [21]))))

	.dataa(\Mux16~10_combout ),
	.datab(\reg_file[11][15]~q ),
	.datac(\reg_file[9][15]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux16~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~11 .lut_mask = 16'hD8AA;
defparam \Mux16~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N16
cycloneive_lcell_comb \Mux16~14 (
// Equation(s):
// \Mux16~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][15]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][15]~q )))))

	.dataa(\reg_file[3][15]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[1][15]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux16~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~14 .lut_mask = 16'hB800;
defparam \Mux16~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N10
cycloneive_lcell_comb \Mux16~15 (
// Equation(s):
// \Mux16~15_combout  = (\Mux16~14_combout ) # ((\prif.imemload_id [22] & (!\prif.imemload_id [21] & \reg_file[2][15]~q )))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\Mux16~14_combout ),
	.datad(\reg_file[2][15]~q ),
	.cin(gnd),
	.combout(\Mux16~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~15 .lut_mask = 16'hF2F0;
defparam \Mux16~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N24
cycloneive_lcell_comb \Mux16~12 (
// Equation(s):
// \Mux16~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][15]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[4][15]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[4][15]~q ),
	.datad(\reg_file[5][15]~q ),
	.cin(gnd),
	.combout(\Mux16~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~12 .lut_mask = 16'hBA98;
defparam \Mux16~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N26
cycloneive_lcell_comb \Mux16~13 (
// Equation(s):
// \Mux16~13_combout  = (\prif.imemload_id [22] & ((\Mux16~12_combout  & ((\reg_file[7][15]~q ))) # (!\Mux16~12_combout  & (\reg_file[6][15]~q )))) # (!\prif.imemload_id [22] & (((\Mux16~12_combout ))))

	.dataa(\reg_file[6][15]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[7][15]~q ),
	.datad(\Mux16~12_combout ),
	.cin(gnd),
	.combout(\Mux16~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~13 .lut_mask = 16'hF388;
defparam \Mux16~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N0
cycloneive_lcell_comb \Mux16~16 (
// Equation(s):
// \Mux16~16_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\Mux16~13_combout ))) # (!\prif.imemload_id [23] & (\Mux16~15_combout ))))

	.dataa(\Mux16~15_combout ),
	.datab(prifimemload_id_24),
	.datac(prifimemload_id_23),
	.datad(\Mux16~13_combout ),
	.cin(gnd),
	.combout(\Mux16~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux16~16 .lut_mask = 16'hF2C2;
defparam \Mux16~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N28
cycloneive_lcell_comb \Mux17~0 (
// Equation(s):
// \Mux17~0_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][14]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][14]~q )))))

	.dataa(\reg_file[25][14]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[17][14]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux17~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~0 .lut_mask = 16'hEE30;
defparam \Mux17~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N4
cycloneive_lcell_comb \Mux17~1 (
// Equation(s):
// \Mux17~1_combout  = (\prif.imemload_id [23] & ((\Mux17~0_combout  & (\reg_file[29][14]~q )) # (!\Mux17~0_combout  & ((\reg_file[21][14]~q ))))) # (!\prif.imemload_id [23] & (((\Mux17~0_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[29][14]~q ),
	.datac(\Mux17~0_combout ),
	.datad(\reg_file[21][14]~q ),
	.cin(gnd),
	.combout(\Mux17~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~1 .lut_mask = 16'hDAD0;
defparam \Mux17~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N0
cycloneive_lcell_comb \Mux17~7 (
// Equation(s):
// \Mux17~7_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[27][14]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[19][14]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][14]~q ),
	.datad(\reg_file[27][14]~q ),
	.cin(gnd),
	.combout(\Mux17~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~7 .lut_mask = 16'hBA98;
defparam \Mux17~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N30
cycloneive_lcell_comb \Mux17~8 (
// Equation(s):
// \Mux17~8_combout  = (\prif.imemload_id [23] & ((\Mux17~7_combout  & (\reg_file[31][14]~q )) # (!\Mux17~7_combout  & ((\reg_file[23][14]~q ))))) # (!\prif.imemload_id [23] & (((\Mux17~7_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[31][14]~q ),
	.datac(\Mux17~7_combout ),
	.datad(\reg_file[23][14]~q ),
	.cin(gnd),
	.combout(\Mux17~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~8 .lut_mask = 16'hDAD0;
defparam \Mux17~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N6
cycloneive_lcell_comb \Mux17~4 (
// Equation(s):
// \Mux17~4_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[20][14]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[16][14]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][14]~q ),
	.datad(\reg_file[20][14]~q ),
	.cin(gnd),
	.combout(\Mux17~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~4 .lut_mask = 16'hBA98;
defparam \Mux17~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N8
cycloneive_lcell_comb \Mux17~5 (
// Equation(s):
// \Mux17~5_combout  = (\prif.imemload_id [24] & ((\Mux17~4_combout  & ((\reg_file[28][14]~q ))) # (!\Mux17~4_combout  & (\reg_file[24][14]~q )))) # (!\prif.imemload_id [24] & (((\Mux17~4_combout ))))

	.dataa(\reg_file[24][14]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[28][14]~q ),
	.datad(\Mux17~4_combout ),
	.cin(gnd),
	.combout(\Mux17~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~5 .lut_mask = 16'hF388;
defparam \Mux17~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N0
cycloneive_lcell_comb \reg_file[30][14]~feeder (
// Equation(s):
// \reg_file[30][14]~feeder_combout  = \reg_file_nxt[31][14]~74_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][14]~74_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[30][14]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[30][14]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[30][14]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N1
dffeas \reg_file[30][14] (
	.clk(!CLK),
	.d(\reg_file[30][14]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][14] .is_wysiwyg = "true";
defparam \reg_file[30][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N16
cycloneive_lcell_comb \Mux17~2 (
// Equation(s):
// \Mux17~2_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[22][14]~q ))) # (!\prif.imemload_id [23] & (\reg_file[18][14]~q ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[18][14]~q ),
	.datac(\reg_file[22][14]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux17~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~2 .lut_mask = 16'hFA44;
defparam \Mux17~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N20
cycloneive_lcell_comb \Mux17~3 (
// Equation(s):
// \Mux17~3_combout  = (\prif.imemload_id [24] & ((\Mux17~2_combout  & (\reg_file[30][14]~q )) # (!\Mux17~2_combout  & ((\reg_file[26][14]~q ))))) # (!\prif.imemload_id [24] & (((\Mux17~2_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[30][14]~q ),
	.datac(\Mux17~2_combout ),
	.datad(\reg_file[26][14]~q ),
	.cin(gnd),
	.combout(\Mux17~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~3 .lut_mask = 16'hDAD0;
defparam \Mux17~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N0
cycloneive_lcell_comb \Mux17~6 (
// Equation(s):
// \Mux17~6_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\Mux17~3_combout ))) # (!\prif.imemload_id [22] & (\Mux17~5_combout ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux17~5_combout ),
	.datad(\Mux17~3_combout ),
	.cin(gnd),
	.combout(\Mux17~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~6 .lut_mask = 16'hDC98;
defparam \Mux17~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N18
cycloneive_lcell_comb \Mux17~15 (
// Equation(s):
// \Mux17~15_combout  = (\Mux17~14_combout ) # ((!\prif.imemload_id [21] & (\prif.imemload_id [22] & \reg_file[2][14]~q )))

	.dataa(\Mux17~14_combout ),
	.datab(prifimemload_id_21),
	.datac(prifimemload_id_22),
	.datad(\reg_file[2][14]~q ),
	.cin(gnd),
	.combout(\Mux17~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~15 .lut_mask = 16'hBAAA;
defparam \Mux17~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N31
dffeas \reg_file[8][14] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][14]~74_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][14]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][14] .is_wysiwyg = "true";
defparam \reg_file[8][14] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N30
cycloneive_lcell_comb \Mux17~12 (
// Equation(s):
// \Mux17~12_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[10][14]~q ))) # (!\prif.imemload_id [22] & (\reg_file[8][14]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[8][14]~q ),
	.datad(\reg_file[10][14]~q ),
	.cin(gnd),
	.combout(\Mux17~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~12 .lut_mask = 16'hDC98;
defparam \Mux17~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N12
cycloneive_lcell_comb \Mux17~13 (
// Equation(s):
// \Mux17~13_combout  = (\Mux17~12_combout  & (((\reg_file[11][14]~q ) # (!\prif.imemload_id [21])))) # (!\Mux17~12_combout  & (\reg_file[9][14]~q  & ((\prif.imemload_id [21]))))

	.dataa(\reg_file[9][14]~q ),
	.datab(\Mux17~12_combout ),
	.datac(\reg_file[11][14]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux17~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~13 .lut_mask = 16'hE2CC;
defparam \Mux17~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N16
cycloneive_lcell_comb \Mux17~16 (
// Equation(s):
// \Mux17~16_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\Mux17~13_combout ))) # (!\prif.imemload_id [24] & (\Mux17~15_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\Mux17~15_combout ),
	.datac(\Mux17~13_combout ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux17~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~16 .lut_mask = 16'hFA44;
defparam \Mux17~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N4
cycloneive_lcell_comb \Mux17~17 (
// Equation(s):
// \Mux17~17_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[13][14]~q ))) # (!\prif.imemload_id [21] & (\reg_file[12][14]~q ))))

	.dataa(\reg_file[12][14]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[13][14]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux17~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~17 .lut_mask = 16'hFC22;
defparam \Mux17~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N6
cycloneive_lcell_comb \Mux17~18 (
// Equation(s):
// \Mux17~18_combout  = (\prif.imemload_id [22] & ((\Mux17~17_combout  & (\reg_file[15][14]~q )) # (!\Mux17~17_combout  & ((\reg_file[14][14]~q ))))) # (!\prif.imemload_id [22] & (((\Mux17~17_combout ))))

	.dataa(\reg_file[15][14]~q ),
	.datab(\reg_file[14][14]~q ),
	.datac(prifimemload_id_22),
	.datad(\Mux17~17_combout ),
	.cin(gnd),
	.combout(\Mux17~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~18 .lut_mask = 16'hAFC0;
defparam \Mux17~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y26_N16
cycloneive_lcell_comb \Mux17~10 (
// Equation(s):
// \Mux17~10_combout  = (\prif.imemload_id [21] & (((\reg_file[5][14]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[4][14]~q  & ((!\prif.imemload_id [22]))))

	.dataa(\reg_file[4][14]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[5][14]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux17~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~10 .lut_mask = 16'hCCE2;
defparam \Mux17~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y27_N24
cycloneive_lcell_comb \Mux17~11 (
// Equation(s):
// \Mux17~11_combout  = (\Mux17~10_combout  & (((\reg_file[7][14]~q ) # (!\prif.imemload_id [22])))) # (!\Mux17~10_combout  & (\reg_file[6][14]~q  & (\prif.imemload_id [22])))

	.dataa(\Mux17~10_combout ),
	.datab(\reg_file[6][14]~q ),
	.datac(prifimemload_id_22),
	.datad(\reg_file[7][14]~q ),
	.cin(gnd),
	.combout(\Mux17~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux17~11 .lut_mask = 16'hEA4A;
defparam \Mux17~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N18
cycloneive_lcell_comb \reg_file[17][13]~feeder (
// Equation(s):
// \reg_file[17][13]~feeder_combout  = \reg_file_nxt[31][13]~75_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][13]~75_combout ),
	.cin(gnd),
	.combout(\reg_file[17][13]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[17][13]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[17][13]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N19
dffeas \reg_file[17][13] (
	.clk(!CLK),
	.d(\reg_file[17][13]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][13] .is_wysiwyg = "true";
defparam \reg_file[17][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N8
cycloneive_lcell_comb \Mux18~0 (
// Equation(s):
// \Mux18~0_combout  = (\prif.imemload_id [23] & ((\reg_file[21][13]~q ) # ((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (((\reg_file[17][13]~q  & !\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[21][13]~q ),
	.datac(\reg_file[17][13]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux18~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~0 .lut_mask = 16'hAAD8;
defparam \Mux18~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N30
cycloneive_lcell_comb \Mux18~1 (
// Equation(s):
// \Mux18~1_combout  = (\prif.imemload_id [24] & ((\Mux18~0_combout  & (\reg_file[29][13]~q )) # (!\Mux18~0_combout  & ((\reg_file[25][13]~q ))))) # (!\prif.imemload_id [24] & (((\Mux18~0_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[29][13]~q ),
	.datac(\Mux18~0_combout ),
	.datad(\reg_file[25][13]~q ),
	.cin(gnd),
	.combout(\Mux18~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~1 .lut_mask = 16'hDAD0;
defparam \Mux18~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N24
cycloneive_lcell_comb \Mux18~7 (
// Equation(s):
// \Mux18~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][13]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][13]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][13]~q ),
	.datad(\reg_file[23][13]~q ),
	.cin(gnd),
	.combout(\Mux18~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~7 .lut_mask = 16'hDC98;
defparam \Mux18~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N20
cycloneive_lcell_comb \Mux18~8 (
// Equation(s):
// \Mux18~8_combout  = (\prif.imemload_id [24] & ((\Mux18~7_combout  & (\reg_file[31][13]~q )) # (!\Mux18~7_combout  & ((\reg_file[27][13]~q ))))) # (!\prif.imemload_id [24] & (\Mux18~7_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux18~7_combout ),
	.datac(\reg_file[31][13]~q ),
	.datad(\reg_file[27][13]~q ),
	.cin(gnd),
	.combout(\Mux18~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~8 .lut_mask = 16'hE6C4;
defparam \Mux18~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y30_N23
dffeas \reg_file[26][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][13] .is_wysiwyg = "true";
defparam \reg_file[26][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N22
cycloneive_lcell_comb \Mux18~2 (
// Equation(s):
// \Mux18~2_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[26][13]~q ))) # (!\prif.imemload_id [24] & (\reg_file[18][13]~q ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[18][13]~q ),
	.datac(\reg_file[26][13]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux18~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~2 .lut_mask = 16'hFA44;
defparam \Mux18~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N14
cycloneive_lcell_comb \Mux18~3 (
// Equation(s):
// \Mux18~3_combout  = (\prif.imemload_id [23] & ((\Mux18~2_combout  & (\reg_file[30][13]~q )) # (!\Mux18~2_combout  & ((\reg_file[22][13]~q ))))) # (!\prif.imemload_id [23] & (\Mux18~2_combout ))

	.dataa(prifimemload_id_23),
	.datab(\Mux18~2_combout ),
	.datac(\reg_file[30][13]~q ),
	.datad(\reg_file[22][13]~q ),
	.cin(gnd),
	.combout(\Mux18~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~3 .lut_mask = 16'hE6C4;
defparam \Mux18~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y34_N13
dffeas \reg_file[28][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][13] .is_wysiwyg = "true";
defparam \reg_file[28][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y34_N27
dffeas \reg_file[16][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][13] .is_wysiwyg = "true";
defparam \reg_file[16][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N26
cycloneive_lcell_comb \Mux18~4 (
// Equation(s):
// \Mux18~4_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[24][13]~q ))) # (!\prif.imemload_id [24] & (\reg_file[16][13]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][13]~q ),
	.datad(\reg_file[24][13]~q ),
	.cin(gnd),
	.combout(\Mux18~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~4 .lut_mask = 16'hDC98;
defparam \Mux18~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N12
cycloneive_lcell_comb \Mux18~5 (
// Equation(s):
// \Mux18~5_combout  = (\prif.imemload_id [23] & ((\Mux18~4_combout  & ((\reg_file[28][13]~q ))) # (!\Mux18~4_combout  & (\reg_file[20][13]~q )))) # (!\prif.imemload_id [23] & (((\Mux18~4_combout ))))

	.dataa(\reg_file[20][13]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[28][13]~q ),
	.datad(\Mux18~4_combout ),
	.cin(gnd),
	.combout(\Mux18~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~5 .lut_mask = 16'hF388;
defparam \Mux18~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N2
cycloneive_lcell_comb \Mux18~6 (
// Equation(s):
// \Mux18~6_combout  = (\prif.imemload_id [22] & ((\Mux18~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((!\prif.imemload_id [21] & \Mux18~5_combout ))))

	.dataa(\Mux18~3_combout ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux18~5_combout ),
	.cin(gnd),
	.combout(\Mux18~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~6 .lut_mask = 16'hCBC8;
defparam \Mux18~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y26_N31
dffeas \reg_file[12][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][13] .is_wysiwyg = "true";
defparam \reg_file[12][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N30
cycloneive_lcell_comb \Mux18~17 (
// Equation(s):
// \Mux18~17_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[13][13]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[12][13]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[12][13]~q ),
	.datad(\reg_file[13][13]~q ),
	.cin(gnd),
	.combout(\Mux18~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~17 .lut_mask = 16'hBA98;
defparam \Mux18~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y24_N8
cycloneive_lcell_comb \Mux18~18 (
// Equation(s):
// \Mux18~18_combout  = (\Mux18~17_combout  & (((\reg_file[15][13]~q ) # (!\prif.imemload_id [22])))) # (!\Mux18~17_combout  & (\reg_file[14][13]~q  & (\prif.imemload_id [22])))

	.dataa(\Mux18~17_combout ),
	.datab(\reg_file[14][13]~q ),
	.datac(prifimemload_id_22),
	.datad(\reg_file[15][13]~q ),
	.cin(gnd),
	.combout(\Mux18~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~18 .lut_mask = 16'hEA4A;
defparam \Mux18~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y35_N27
dffeas \reg_file[8][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][13] .is_wysiwyg = "true";
defparam \reg_file[8][13] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y35_N13
dffeas \reg_file[10][13] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][13]~75_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][13]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][13] .is_wysiwyg = "true";
defparam \reg_file[10][13] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y35_N26
cycloneive_lcell_comb \Mux18~10 (
// Equation(s):
// \Mux18~10_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[10][13]~q ))) # (!\prif.imemload_id [22] & (\reg_file[8][13]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[8][13]~q ),
	.datad(\reg_file[10][13]~q ),
	.cin(gnd),
	.combout(\Mux18~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~10 .lut_mask = 16'hDC98;
defparam \Mux18~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N20
cycloneive_lcell_comb \Mux18~11 (
// Equation(s):
// \Mux18~11_combout  = (\Mux18~10_combout  & (((\reg_file[11][13]~q )) # (!\prif.imemload_id [21]))) # (!\Mux18~10_combout  & (\prif.imemload_id [21] & (\reg_file[9][13]~q )))

	.dataa(\Mux18~10_combout ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[9][13]~q ),
	.datad(\reg_file[11][13]~q ),
	.cin(gnd),
	.combout(\Mux18~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~11 .lut_mask = 16'hEA62;
defparam \Mux18~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N4
cycloneive_lcell_comb \Mux18~14 (
// Equation(s):
// \Mux18~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][13]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][13]~q ))))

	.dataa(\reg_file[1][13]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][13]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux18~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~14 .lut_mask = 16'hE200;
defparam \Mux18~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N14
cycloneive_lcell_comb \Mux18~15 (
// Equation(s):
// \Mux18~15_combout  = (\Mux18~14_combout ) # ((\reg_file[2][13]~q  & (\prif.imemload_id [22] & !\prif.imemload_id [21])))

	.dataa(\reg_file[2][13]~q ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux18~14_combout ),
	.cin(gnd),
	.combout(\Mux18~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~15 .lut_mask = 16'hFF08;
defparam \Mux18~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N18
cycloneive_lcell_comb \Mux18~13 (
// Equation(s):
// \Mux18~13_combout  = (\Mux18~12_combout  & (((\reg_file[7][13]~q )) # (!\prif.imemload_id [22]))) # (!\Mux18~12_combout  & (\prif.imemload_id [22] & ((\reg_file[6][13]~q ))))

	.dataa(\Mux18~12_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[7][13]~q ),
	.datad(\reg_file[6][13]~q ),
	.cin(gnd),
	.combout(\Mux18~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~13 .lut_mask = 16'hE6A2;
defparam \Mux18~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y24_N0
cycloneive_lcell_comb \Mux18~16 (
// Equation(s):
// \Mux18~16_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\Mux18~13_combout ))) # (!\prif.imemload_id [23] & (\Mux18~15_combout ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\Mux18~15_combout ),
	.datad(\Mux18~13_combout ),
	.cin(gnd),
	.combout(\Mux18~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux18~16 .lut_mask = 16'hDC98;
defparam \Mux18~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y30_N30
cycloneive_lcell_comb \Mux20~2 (
// Equation(s):
// \Mux20~2_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[26][11]~q ))) # (!\prif.imemload_id [24] & (\reg_file[18][11]~q ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[18][11]~q ),
	.datac(\reg_file[26][11]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux20~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~2 .lut_mask = 16'hFA44;
defparam \Mux20~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N2
cycloneive_lcell_comb \Mux20~3 (
// Equation(s):
// \Mux20~3_combout  = (\prif.imemload_id [23] & ((\Mux20~2_combout  & ((\reg_file[30][11]~q ))) # (!\Mux20~2_combout  & (\reg_file[22][11]~q )))) # (!\prif.imemload_id [23] & (((\Mux20~2_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[22][11]~q ),
	.datac(\reg_file[30][11]~q ),
	.datad(\Mux20~2_combout ),
	.cin(gnd),
	.combout(\Mux20~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~3 .lut_mask = 16'hF588;
defparam \Mux20~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y34_N14
cycloneive_lcell_comb \Mux20~4 (
// Equation(s):
// \Mux20~4_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[24][11]~q ))) # (!\prif.imemload_id [24] & (\reg_file[16][11]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][11]~q ),
	.datad(\reg_file[24][11]~q ),
	.cin(gnd),
	.combout(\Mux20~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~4 .lut_mask = 16'hDC98;
defparam \Mux20~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N8
cycloneive_lcell_comb \Mux20~5 (
// Equation(s):
// \Mux20~5_combout  = (\Mux20~4_combout  & (((\reg_file[28][11]~q ) # (!\prif.imemload_id [23])))) # (!\Mux20~4_combout  & (\reg_file[20][11]~q  & ((\prif.imemload_id [23]))))

	.dataa(\reg_file[20][11]~q ),
	.datab(\Mux20~4_combout ),
	.datac(\reg_file[28][11]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux20~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~5 .lut_mask = 16'hE2CC;
defparam \Mux20~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N20
cycloneive_lcell_comb \Mux20~6 (
// Equation(s):
// \Mux20~6_combout  = (\prif.imemload_id [22] & ((\Mux20~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((!\prif.imemload_id [21] & \Mux20~5_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\Mux20~3_combout ),
	.datac(prifimemload_id_21),
	.datad(\Mux20~5_combout ),
	.cin(gnd),
	.combout(\Mux20~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~6 .lut_mask = 16'hADA8;
defparam \Mux20~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N31
dffeas \reg_file[17][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][11] .is_wysiwyg = "true";
defparam \reg_file[17][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N30
cycloneive_lcell_comb \Mux20~0 (
// Equation(s):
// \Mux20~0_combout  = (\prif.imemload_id [23] & ((\reg_file[21][11]~q ) # ((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (((\reg_file[17][11]~q  & !\prif.imemload_id [24]))))

	.dataa(\reg_file[21][11]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[17][11]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux20~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~0 .lut_mask = 16'hCCB8;
defparam \Mux20~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N10
cycloneive_lcell_comb \Mux20~1 (
// Equation(s):
// \Mux20~1_combout  = (\prif.imemload_id [24] & ((\Mux20~0_combout  & (\reg_file[29][11]~q )) # (!\Mux20~0_combout  & ((\reg_file[25][11]~q ))))) # (!\prif.imemload_id [24] & (\Mux20~0_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux20~0_combout ),
	.datac(\reg_file[29][11]~q ),
	.datad(\reg_file[25][11]~q ),
	.cin(gnd),
	.combout(\Mux20~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~1 .lut_mask = 16'hE6C4;
defparam \Mux20~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N28
cycloneive_lcell_comb \Mux20~7 (
// Equation(s):
// \Mux20~7_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\reg_file[23][11]~q )) # (!\prif.imemload_id [23] & ((\reg_file[19][11]~q )))))

	.dataa(\reg_file[23][11]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[19][11]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux20~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~7 .lut_mask = 16'hEE30;
defparam \Mux20~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N10
cycloneive_lcell_comb \Mux20~8 (
// Equation(s):
// \Mux20~8_combout  = (\prif.imemload_id [24] & ((\Mux20~7_combout  & (\reg_file[31][11]~q )) # (!\Mux20~7_combout  & ((\reg_file[27][11]~q ))))) # (!\prif.imemload_id [24] & (((\Mux20~7_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[31][11]~q ),
	.datac(\reg_file[27][11]~q ),
	.datad(\Mux20~7_combout ),
	.cin(gnd),
	.combout(\Mux20~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~8 .lut_mask = 16'hDDA0;
defparam \Mux20~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N28
cycloneive_lcell_comb \Mux20~12 (
// Equation(s):
// \Mux20~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][11]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[4][11]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[4][11]~q ),
	.datad(\reg_file[5][11]~q ),
	.cin(gnd),
	.combout(\Mux20~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~12 .lut_mask = 16'hBA98;
defparam \Mux20~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N6
cycloneive_lcell_comb \Mux20~13 (
// Equation(s):
// \Mux20~13_combout  = (\prif.imemload_id [22] & ((\Mux20~12_combout  & ((\reg_file[7][11]~q ))) # (!\Mux20~12_combout  & (\reg_file[6][11]~q )))) # (!\prif.imemload_id [22] & (((\Mux20~12_combout ))))

	.dataa(\reg_file[6][11]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[7][11]~q ),
	.datad(\Mux20~12_combout ),
	.cin(gnd),
	.combout(\Mux20~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~13 .lut_mask = 16'hF388;
defparam \Mux20~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N14
cycloneive_lcell_comb \Mux20~14 (
// Equation(s):
// \Mux20~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][11]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][11]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[1][11]~q ),
	.datad(\reg_file[3][11]~q ),
	.cin(gnd),
	.combout(\Mux20~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~14 .lut_mask = 16'hA820;
defparam \Mux20~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N30
cycloneive_lcell_comb \Mux20~15 (
// Equation(s):
// \Mux20~15_combout  = (\Mux20~14_combout ) # ((!\prif.imemload_id [21] & (\prif.imemload_id [22] & \reg_file[2][11]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux20~14_combout ),
	.datad(\reg_file[2][11]~q ),
	.cin(gnd),
	.combout(\Mux20~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~15 .lut_mask = 16'hF4F0;
defparam \Mux20~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N18
cycloneive_lcell_comb \Mux20~16 (
// Equation(s):
// \Mux20~16_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\Mux20~13_combout )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & ((\Mux20~15_combout ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux20~13_combout ),
	.datad(\Mux20~15_combout ),
	.cin(gnd),
	.combout(\Mux20~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~16 .lut_mask = 16'hB9A8;
defparam \Mux20~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N7
dffeas \reg_file[8][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][11] .is_wysiwyg = "true";
defparam \reg_file[8][11] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N17
dffeas \reg_file[10][11] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][11]~77_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][11]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][11] .is_wysiwyg = "true";
defparam \reg_file[10][11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N6
cycloneive_lcell_comb \Mux20~10 (
// Equation(s):
// \Mux20~10_combout  = (\prif.imemload_id [22] & ((\prif.imemload_id [21]) # ((\reg_file[10][11]~q )))) # (!\prif.imemload_id [22] & (!\prif.imemload_id [21] & (\reg_file[8][11]~q )))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[8][11]~q ),
	.datad(\reg_file[10][11]~q ),
	.cin(gnd),
	.combout(\Mux20~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~10 .lut_mask = 16'hBA98;
defparam \Mux20~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N24
cycloneive_lcell_comb \Mux20~11 (
// Equation(s):
// \Mux20~11_combout  = (\Mux20~10_combout  & ((\reg_file[11][11]~q ) # ((!\prif.imemload_id [21])))) # (!\Mux20~10_combout  & (((\reg_file[9][11]~q  & \prif.imemload_id [21]))))

	.dataa(\reg_file[11][11]~q ),
	.datab(\Mux20~10_combout ),
	.datac(\reg_file[9][11]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux20~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~11 .lut_mask = 16'hB8CC;
defparam \Mux20~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N18
cycloneive_lcell_comb \Mux20~17 (
// Equation(s):
// \Mux20~17_combout  = (\prif.imemload_id [21] & ((\reg_file[13][11]~q ) # ((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (((\reg_file[12][11]~q  & !\prif.imemload_id [22]))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[13][11]~q ),
	.datac(\reg_file[12][11]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux20~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~17 .lut_mask = 16'hAAD8;
defparam \Mux20~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N0
cycloneive_lcell_comb \Mux20~18 (
// Equation(s):
// \Mux20~18_combout  = (\prif.imemload_id [22] & ((\Mux20~17_combout  & ((\reg_file[15][11]~q ))) # (!\Mux20~17_combout  & (\reg_file[14][11]~q )))) # (!\prif.imemload_id [22] & (((\Mux20~17_combout ))))

	.dataa(\reg_file[14][11]~q ),
	.datab(prifimemload_id_22),
	.datac(\Mux20~17_combout ),
	.datad(\reg_file[15][11]~q ),
	.cin(gnd),
	.combout(\Mux20~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux20~18 .lut_mask = 16'hF838;
defparam \Mux20~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N4
cycloneive_lcell_comb \Mux19~7 (
// Equation(s):
// \Mux19~7_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[27][12]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[19][12]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][12]~q ),
	.datad(\reg_file[27][12]~q ),
	.cin(gnd),
	.combout(\Mux19~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~7 .lut_mask = 16'hBA98;
defparam \Mux19~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y26_N30
cycloneive_lcell_comb \Mux19~8 (
// Equation(s):
// \Mux19~8_combout  = (\prif.imemload_id [23] & ((\Mux19~7_combout  & ((\reg_file[31][12]~q ))) # (!\Mux19~7_combout  & (\reg_file[23][12]~q )))) # (!\prif.imemload_id [23] & (((\Mux19~7_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[23][12]~q ),
	.datac(\reg_file[31][12]~q ),
	.datad(\Mux19~7_combout ),
	.cin(gnd),
	.combout(\Mux19~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~8 .lut_mask = 16'hF588;
defparam \Mux19~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N24
cycloneive_lcell_comb \Mux19~0 (
// Equation(s):
// \Mux19~0_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][12]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][12]~q )))))

	.dataa(\reg_file[25][12]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[17][12]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux19~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~0 .lut_mask = 16'hEE30;
defparam \Mux19~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N6
cycloneive_lcell_comb \Mux19~1 (
// Equation(s):
// \Mux19~1_combout  = (\prif.imemload_id [23] & ((\Mux19~0_combout  & (\reg_file[29][12]~q )) # (!\Mux19~0_combout  & ((\reg_file[21][12]~q ))))) # (!\prif.imemload_id [23] & (((\Mux19~0_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[29][12]~q ),
	.datac(\Mux19~0_combout ),
	.datad(\reg_file[21][12]~q ),
	.cin(gnd),
	.combout(\Mux19~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~1 .lut_mask = 16'hDAD0;
defparam \Mux19~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N8
cycloneive_lcell_comb \Mux19~3 (
// Equation(s):
// \Mux19~3_combout  = (\Mux19~2_combout  & (((\reg_file[30][12]~q ) # (!\prif.imemload_id [24])))) # (!\Mux19~2_combout  & (\reg_file[26][12]~q  & ((\prif.imemload_id [24]))))

	.dataa(\Mux19~2_combout ),
	.datab(\reg_file[26][12]~q ),
	.datac(\reg_file[30][12]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux19~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~3 .lut_mask = 16'hE4AA;
defparam \Mux19~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N20
cycloneive_lcell_comb \Mux19~4 (
// Equation(s):
// \Mux19~4_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\reg_file[20][12]~q )) # (!\prif.imemload_id [23] & ((\reg_file[16][12]~q )))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[20][12]~q ),
	.datac(\reg_file[16][12]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux19~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~4 .lut_mask = 16'hEE50;
defparam \Mux19~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N2
cycloneive_lcell_comb \Mux19~5 (
// Equation(s):
// \Mux19~5_combout  = (\prif.imemload_id [24] & ((\Mux19~4_combout  & (\reg_file[28][12]~q )) # (!\Mux19~4_combout  & ((\reg_file[24][12]~q ))))) # (!\prif.imemload_id [24] & (((\Mux19~4_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[28][12]~q ),
	.datac(\reg_file[24][12]~q ),
	.datad(\Mux19~4_combout ),
	.cin(gnd),
	.combout(\Mux19~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~5 .lut_mask = 16'hDDA0;
defparam \Mux19~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N6
cycloneive_lcell_comb \Mux19~6 (
// Equation(s):
// \Mux19~6_combout  = (\prif.imemload_id [22] & ((\Mux19~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((!\prif.imemload_id [21] & \Mux19~5_combout ))))

	.dataa(\Mux19~3_combout ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux19~5_combout ),
	.cin(gnd),
	.combout(\Mux19~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~6 .lut_mask = 16'hCBC8;
defparam \Mux19~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y26_N26
cycloneive_lcell_comb \reg_file[6][12]~feeder (
// Equation(s):
// \reg_file[6][12]~feeder_combout  = \reg_file_nxt[31][12]~76_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][12]~76_combout ),
	.cin(gnd),
	.combout(\reg_file[6][12]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][12]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[6][12]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y26_N27
dffeas \reg_file[6][12] (
	.clk(!CLK),
	.d(\reg_file[6][12]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][12]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][12] .is_wysiwyg = "true";
defparam \reg_file[6][12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N20
cycloneive_lcell_comb \Mux19~10 (
// Equation(s):
// \Mux19~10_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[5][12]~q ))) # (!\prif.imemload_id [21] & (\reg_file[4][12]~q ))))

	.dataa(\reg_file[4][12]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[5][12]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux19~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~10 .lut_mask = 16'hFC22;
defparam \Mux19~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y27_N8
cycloneive_lcell_comb \Mux19~11 (
// Equation(s):
// \Mux19~11_combout  = (\prif.imemload_id [22] & ((\Mux19~10_combout  & ((\reg_file[7][12]~q ))) # (!\Mux19~10_combout  & (\reg_file[6][12]~q )))) # (!\prif.imemload_id [22] & (((\Mux19~10_combout ))))

	.dataa(\reg_file[6][12]~q ),
	.datab(\reg_file[7][12]~q ),
	.datac(prifimemload_id_22),
	.datad(\Mux19~10_combout ),
	.cin(gnd),
	.combout(\Mux19~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~11 .lut_mask = 16'hCFA0;
defparam \Mux19~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N0
cycloneive_lcell_comb \Mux19~17 (
// Equation(s):
// \Mux19~17_combout  = (\prif.imemload_id [21] & (((\reg_file[13][12]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[12][12]~q  & ((!\prif.imemload_id [22]))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[12][12]~q ),
	.datac(\reg_file[13][12]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux19~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~17 .lut_mask = 16'hAAE4;
defparam \Mux19~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N10
cycloneive_lcell_comb \Mux19~18 (
// Equation(s):
// \Mux19~18_combout  = (\prif.imemload_id [22] & ((\Mux19~17_combout  & ((\reg_file[15][12]~q ))) # (!\Mux19~17_combout  & (\reg_file[14][12]~q )))) # (!\prif.imemload_id [22] & (((\Mux19~17_combout ))))

	.dataa(\reg_file[14][12]~q ),
	.datab(prifimemload_id_22),
	.datac(\Mux19~17_combout ),
	.datad(\reg_file[15][12]~q ),
	.cin(gnd),
	.combout(\Mux19~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~18 .lut_mask = 16'hF838;
defparam \Mux19~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N22
cycloneive_lcell_comb \Mux19~13 (
// Equation(s):
// \Mux19~13_combout  = (\Mux19~12_combout  & (((\reg_file[11][12]~q ) # (!\prif.imemload_id [21])))) # (!\Mux19~12_combout  & (\reg_file[9][12]~q  & ((\prif.imemload_id [21]))))

	.dataa(\Mux19~12_combout ),
	.datab(\reg_file[9][12]~q ),
	.datac(\reg_file[11][12]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux19~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~13 .lut_mask = 16'hE4AA;
defparam \Mux19~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N22
cycloneive_lcell_comb \Mux19~15 (
// Equation(s):
// \Mux19~15_combout  = (\Mux19~14_combout ) # ((\reg_file[2][12]~q  & (!\prif.imemload_id [21] & \prif.imemload_id [22])))

	.dataa(\Mux19~14_combout ),
	.datab(\reg_file[2][12]~q ),
	.datac(prifimemload_id_21),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux19~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~15 .lut_mask = 16'hAEAA;
defparam \Mux19~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N16
cycloneive_lcell_comb \Mux19~16 (
// Equation(s):
// \Mux19~16_combout  = (\prif.imemload_id [24] & ((\Mux19~13_combout ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\Mux19~15_combout  & !\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\Mux19~13_combout ),
	.datac(\Mux19~15_combout ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux19~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux19~16 .lut_mask = 16'hAAD8;
defparam \Mux19~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N20
cycloneive_lcell_comb \Mux21~7 (
// Equation(s):
// \Mux21~7_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[27][10]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[19][10]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][10]~q ),
	.datad(\reg_file[27][10]~q ),
	.cin(gnd),
	.combout(\Mux21~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~7 .lut_mask = 16'hBA98;
defparam \Mux21~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N12
cycloneive_lcell_comb \Mux21~8 (
// Equation(s):
// \Mux21~8_combout  = (\Mux21~7_combout  & (((\reg_file[31][10]~q ) # (!\prif.imemload_id [23])))) # (!\Mux21~7_combout  & (\reg_file[23][10]~q  & ((\prif.imemload_id [23]))))

	.dataa(\Mux21~7_combout ),
	.datab(\reg_file[23][10]~q ),
	.datac(\reg_file[31][10]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux21~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~8 .lut_mask = 16'hE4AA;
defparam \Mux21~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y30_N18
cycloneive_lcell_comb \Mux21~2 (
// Equation(s):
// \Mux21~2_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[22][10]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & ((\reg_file[18][10]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[22][10]~q ),
	.datad(\reg_file[18][10]~q ),
	.cin(gnd),
	.combout(\Mux21~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~2 .lut_mask = 16'hB9A8;
defparam \Mux21~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N2
cycloneive_lcell_comb \Mux21~3 (
// Equation(s):
// \Mux21~3_combout  = (\prif.imemload_id [24] & ((\Mux21~2_combout  & (\reg_file[30][10]~q )) # (!\Mux21~2_combout  & ((\reg_file[26][10]~q ))))) # (!\prif.imemload_id [24] & (((\Mux21~2_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[30][10]~q ),
	.datac(\reg_file[26][10]~q ),
	.datad(\Mux21~2_combout ),
	.cin(gnd),
	.combout(\Mux21~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~3 .lut_mask = 16'hDDA0;
defparam \Mux21~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N4
cycloneive_lcell_comb \Mux21~4 (
// Equation(s):
// \Mux21~4_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[20][10]~q ))) # (!\prif.imemload_id [23] & (\reg_file[16][10]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[16][10]~q ),
	.datad(\reg_file[20][10]~q ),
	.cin(gnd),
	.combout(\Mux21~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~4 .lut_mask = 16'hDC98;
defparam \Mux21~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N31
dffeas \reg_file[28][10] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][10]~78_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~29_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[28][10]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[28][10] .is_wysiwyg = "true";
defparam \reg_file[28][10] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N30
cycloneive_lcell_comb \Mux21~5 (
// Equation(s):
// \Mux21~5_combout  = (\prif.imemload_id [24] & ((\Mux21~4_combout  & (\reg_file[28][10]~q )) # (!\Mux21~4_combout  & ((\reg_file[24][10]~q ))))) # (!\prif.imemload_id [24] & (\Mux21~4_combout ))

	.dataa(prifimemload_id_24),
	.datab(\Mux21~4_combout ),
	.datac(\reg_file[28][10]~q ),
	.datad(\reg_file[24][10]~q ),
	.cin(gnd),
	.combout(\Mux21~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~5 .lut_mask = 16'hE6C4;
defparam \Mux21~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N18
cycloneive_lcell_comb \Mux21~6 (
// Equation(s):
// \Mux21~6_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\Mux21~3_combout )) # (!\prif.imemload_id [22] & ((\Mux21~5_combout )))))

	.dataa(\Mux21~3_combout ),
	.datab(prifimemload_id_21),
	.datac(prifimemload_id_22),
	.datad(\Mux21~5_combout ),
	.cin(gnd),
	.combout(\Mux21~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~6 .lut_mask = 16'hE3E0;
defparam \Mux21~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N8
cycloneive_lcell_comb \Mux21~0 (
// Equation(s):
// \Mux21~0_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][10]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][10]~q )))))

	.dataa(\reg_file[25][10]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[17][10]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux21~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~0 .lut_mask = 16'hEE30;
defparam \Mux21~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y28_N20
cycloneive_lcell_comb \Mux21~1 (
// Equation(s):
// \Mux21~1_combout  = (\prif.imemload_id [23] & ((\Mux21~0_combout  & (\reg_file[29][10]~q )) # (!\Mux21~0_combout  & ((\reg_file[21][10]~q ))))) # (!\prif.imemload_id [23] & (\Mux21~0_combout ))

	.dataa(prifimemload_id_23),
	.datab(\Mux21~0_combout ),
	.datac(\reg_file[29][10]~q ),
	.datad(\reg_file[21][10]~q ),
	.cin(gnd),
	.combout(\Mux21~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~1 .lut_mask = 16'hE6C4;
defparam \Mux21~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N2
cycloneive_lcell_comb \Mux21~10 (
// Equation(s):
// \Mux21~10_combout  = (\prif.imemload_id [21] & ((\reg_file[5][10]~q ) # ((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (((\reg_file[4][10]~q  & !\prif.imemload_id [22]))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[5][10]~q ),
	.datac(\reg_file[4][10]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux21~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~10 .lut_mask = 16'hAAD8;
defparam \Mux21~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N24
cycloneive_lcell_comb \Mux21~11 (
// Equation(s):
// \Mux21~11_combout  = (\prif.imemload_id [22] & ((\Mux21~10_combout  & ((\reg_file[7][10]~q ))) # (!\Mux21~10_combout  & (\reg_file[6][10]~q )))) # (!\prif.imemload_id [22] & (\Mux21~10_combout ))

	.dataa(prifimemload_id_22),
	.datab(\Mux21~10_combout ),
	.datac(\reg_file[6][10]~q ),
	.datad(\reg_file[7][10]~q ),
	.cin(gnd),
	.combout(\Mux21~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~11 .lut_mask = 16'hEC64;
defparam \Mux21~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N16
cycloneive_lcell_comb \Mux21~17 (
// Equation(s):
// \Mux21~17_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[13][10]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & ((\reg_file[12][10]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[13][10]~q ),
	.datad(\reg_file[12][10]~q ),
	.cin(gnd),
	.combout(\Mux21~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~17 .lut_mask = 16'hB9A8;
defparam \Mux21~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N18
cycloneive_lcell_comb \Mux21~18 (
// Equation(s):
// \Mux21~18_combout  = (\Mux21~17_combout  & ((\reg_file[15][10]~q ) # ((!\prif.imemload_id [22])))) # (!\Mux21~17_combout  & (((\prif.imemload_id [22] & \reg_file[14][10]~q ))))

	.dataa(\Mux21~17_combout ),
	.datab(\reg_file[15][10]~q ),
	.datac(prifimemload_id_22),
	.datad(\reg_file[14][10]~q ),
	.cin(gnd),
	.combout(\Mux21~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~18 .lut_mask = 16'hDA8A;
defparam \Mux21~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N0
cycloneive_lcell_comb \Mux21~14 (
// Equation(s):
// \Mux21~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][10]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][10]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[1][10]~q ),
	.datad(\reg_file[3][10]~q ),
	.cin(gnd),
	.combout(\Mux21~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~14 .lut_mask = 16'hA820;
defparam \Mux21~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N30
cycloneive_lcell_comb \Mux21~15 (
// Equation(s):
// \Mux21~15_combout  = (\Mux21~14_combout ) # ((!\prif.imemload_id [21] & (\reg_file[2][10]~q  & \prif.imemload_id [22])))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[2][10]~q ),
	.datac(\Mux21~14_combout ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux21~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~15 .lut_mask = 16'hF4F0;
defparam \Mux21~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N2
cycloneive_lcell_comb \Mux21~13 (
// Equation(s):
// \Mux21~13_combout  = (\Mux21~12_combout  & (((\reg_file[11][10]~q )) # (!\prif.imemload_id [21]))) # (!\Mux21~12_combout  & (\prif.imemload_id [21] & ((\reg_file[9][10]~q ))))

	.dataa(\Mux21~12_combout ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[11][10]~q ),
	.datad(\reg_file[9][10]~q ),
	.cin(gnd),
	.combout(\Mux21~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~13 .lut_mask = 16'hE6A2;
defparam \Mux21~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y25_N20
cycloneive_lcell_comb \Mux21~16 (
// Equation(s):
// \Mux21~16_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\Mux21~13_combout ))) # (!\prif.imemload_id [24] & (\Mux21~15_combout ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux21~15_combout ),
	.datad(\Mux21~13_combout ),
	.cin(gnd),
	.combout(\Mux21~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux21~16 .lut_mask = 16'hDC98;
defparam \Mux21~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N22
cycloneive_lcell_comb \Mux22~0 (
// Equation(s):
// \Mux22~0_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[21][9]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[17][9]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[17][9]~q ),
	.datad(\reg_file[21][9]~q ),
	.cin(gnd),
	.combout(\Mux22~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~0 .lut_mask = 16'hBA98;
defparam \Mux22~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N8
cycloneive_lcell_comb \Mux22~1 (
// Equation(s):
// \Mux22~1_combout  = (\Mux22~0_combout  & (((\reg_file[29][9]~q ) # (!\prif.imemload_id [24])))) # (!\Mux22~0_combout  & (\reg_file[25][9]~q  & ((\prif.imemload_id [24]))))

	.dataa(\Mux22~0_combout ),
	.datab(\reg_file[25][9]~q ),
	.datac(\reg_file[29][9]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux22~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~1 .lut_mask = 16'hE4AA;
defparam \Mux22~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N7
dffeas \reg_file[19][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][9] .is_wysiwyg = "true";
defparam \reg_file[19][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N6
cycloneive_lcell_comb \Mux22~7 (
// Equation(s):
// \Mux22~7_combout  = (\prif.imemload_id [23] & ((\reg_file[23][9]~q ) # ((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (((\reg_file[19][9]~q  & !\prif.imemload_id [24]))))

	.dataa(\reg_file[23][9]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][9]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux22~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~7 .lut_mask = 16'hCCB8;
defparam \Mux22~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N8
cycloneive_lcell_comb \Mux22~8 (
// Equation(s):
// \Mux22~8_combout  = (\Mux22~7_combout  & (((\reg_file[31][9]~q )) # (!\prif.imemload_id [24]))) # (!\Mux22~7_combout  & (\prif.imemload_id [24] & ((\reg_file[27][9]~q ))))

	.dataa(\Mux22~7_combout ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[31][9]~q ),
	.datad(\reg_file[27][9]~q ),
	.cin(gnd),
	.combout(\Mux22~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~8 .lut_mask = 16'hE6A2;
defparam \Mux22~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N12
cycloneive_lcell_comb \Mux22~4 (
// Equation(s):
// \Mux22~4_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[24][9]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & ((\reg_file[16][9]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[24][9]~q ),
	.datad(\reg_file[16][9]~q ),
	.cin(gnd),
	.combout(\Mux22~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~4 .lut_mask = 16'hB9A8;
defparam \Mux22~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N2
cycloneive_lcell_comb \Mux22~5 (
// Equation(s):
// \Mux22~5_combout  = (\prif.imemload_id [23] & ((\Mux22~4_combout  & ((\reg_file[28][9]~q ))) # (!\Mux22~4_combout  & (\reg_file[20][9]~q )))) # (!\prif.imemload_id [23] & (((\Mux22~4_combout ))))

	.dataa(\reg_file[20][9]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[28][9]~q ),
	.datad(\Mux22~4_combout ),
	.cin(gnd),
	.combout(\Mux22~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~5 .lut_mask = 16'hF388;
defparam \Mux22~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y29_N0
cycloneive_lcell_comb \Mux22~3 (
// Equation(s):
// \Mux22~3_combout  = (\Mux22~2_combout  & (((\reg_file[30][9]~q )) # (!\prif.imemload_id [23]))) # (!\Mux22~2_combout  & (\prif.imemload_id [23] & (\reg_file[22][9]~q )))

	.dataa(\Mux22~2_combout ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[22][9]~q ),
	.datad(\reg_file[30][9]~q ),
	.cin(gnd),
	.combout(\Mux22~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~3 .lut_mask = 16'hEA62;
defparam \Mux22~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N4
cycloneive_lcell_comb \Mux22~6 (
// Equation(s):
// \Mux22~6_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\Mux22~3_combout ))) # (!\prif.imemload_id [22] & (\Mux22~5_combout ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux22~5_combout ),
	.datad(\Mux22~3_combout ),
	.cin(gnd),
	.combout(\Mux22~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~6 .lut_mask = 16'hDC98;
defparam \Mux22~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N0
cycloneive_lcell_comb \Mux22~17 (
// Equation(s):
// \Mux22~17_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[13][9]~q ))) # (!\prif.imemload_id [21] & (\reg_file[12][9]~q ))))

	.dataa(\reg_file[12][9]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[13][9]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux22~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~17 .lut_mask = 16'hFC22;
defparam \Mux22~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y31_N4
cycloneive_lcell_comb \Mux22~18 (
// Equation(s):
// \Mux22~18_combout  = (\Mux22~17_combout  & (((\reg_file[15][9]~q )) # (!\prif.imemload_id [22]))) # (!\Mux22~17_combout  & (\prif.imemload_id [22] & (\reg_file[14][9]~q )))

	.dataa(\Mux22~17_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[14][9]~q ),
	.datad(\reg_file[15][9]~q ),
	.cin(gnd),
	.combout(\Mux22~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~18 .lut_mask = 16'hEA62;
defparam \Mux22~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y33_N29
dffeas \reg_file[10][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~35_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[10][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[10][9] .is_wysiwyg = "true";
defparam \reg_file[10][9] .power_up = "low";
// synopsys translate_on

// Location: FF_X69_Y33_N11
dffeas \reg_file[8][9] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][9]~79_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][9]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][9] .is_wysiwyg = "true";
defparam \reg_file[8][9] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N28
cycloneive_lcell_comb \Mux22~10 (
// Equation(s):
// \Mux22~10_combout  = (\prif.imemload_id [22] & ((\prif.imemload_id [21]) # ((\reg_file[10][9]~q )))) # (!\prif.imemload_id [22] & (!\prif.imemload_id [21] & ((\reg_file[8][9]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[10][9]~q ),
	.datad(\reg_file[8][9]~q ),
	.cin(gnd),
	.combout(\Mux22~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~10 .lut_mask = 16'hB9A8;
defparam \Mux22~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y31_N8
cycloneive_lcell_comb \Mux22~11 (
// Equation(s):
// \Mux22~11_combout  = (\prif.imemload_id [21] & ((\Mux22~10_combout  & ((\reg_file[11][9]~q ))) # (!\Mux22~10_combout  & (\reg_file[9][9]~q )))) # (!\prif.imemload_id [21] & (\Mux22~10_combout ))

	.dataa(prifimemload_id_21),
	.datab(\Mux22~10_combout ),
	.datac(\reg_file[9][9]~q ),
	.datad(\reg_file[11][9]~q ),
	.cin(gnd),
	.combout(\Mux22~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~11 .lut_mask = 16'hEC64;
defparam \Mux22~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N8
cycloneive_lcell_comb \Mux22~15 (
// Equation(s):
// \Mux22~15_combout  = (\Mux22~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][9]~q  & !\prif.imemload_id [21])))

	.dataa(\Mux22~14_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][9]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux22~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~15 .lut_mask = 16'hAAEA;
defparam \Mux22~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N20
cycloneive_lcell_comb \Mux22~12 (
// Equation(s):
// \Mux22~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][9]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[4][9]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[4][9]~q ),
	.datad(\reg_file[5][9]~q ),
	.cin(gnd),
	.combout(\Mux22~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~12 .lut_mask = 16'hBA98;
defparam \Mux22~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N2
cycloneive_lcell_comb \Mux22~13 (
// Equation(s):
// \Mux22~13_combout  = (\prif.imemload_id [22] & ((\Mux22~12_combout  & ((\reg_file[7][9]~q ))) # (!\Mux22~12_combout  & (\reg_file[6][9]~q )))) # (!\prif.imemload_id [22] & (((\Mux22~12_combout ))))

	.dataa(\reg_file[6][9]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[7][9]~q ),
	.datad(\Mux22~12_combout ),
	.cin(gnd),
	.combout(\Mux22~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~13 .lut_mask = 16'hF388;
defparam \Mux22~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y25_N6
cycloneive_lcell_comb \Mux22~16 (
// Equation(s):
// \Mux22~16_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24]) # (\Mux22~13_combout )))) # (!\prif.imemload_id [23] & (\Mux22~15_combout  & (!\prif.imemload_id [24])))

	.dataa(prifimemload_id_23),
	.datab(\Mux22~15_combout ),
	.datac(prifimemload_id_24),
	.datad(\Mux22~13_combout ),
	.cin(gnd),
	.combout(\Mux22~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux22~16 .lut_mask = 16'hAEA4;
defparam \Mux22~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N8
cycloneive_lcell_comb \Mux13~7 (
// Equation(s):
// \Mux13~7_combout  = (\prif.imemload_id [24] & ((\reg_file[27][18]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[19][18]~q  & !\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[27][18]~q ),
	.datac(\reg_file[19][18]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux13~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~7 .lut_mask = 16'hAAD8;
defparam \Mux13~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N14
cycloneive_lcell_comb \Mux13~8 (
// Equation(s):
// \Mux13~8_combout  = (\Mux13~7_combout  & (((\reg_file[31][18]~q ) # (!\prif.imemload_id [23])))) # (!\Mux13~7_combout  & (\reg_file[23][18]~q  & ((\prif.imemload_id [23]))))

	.dataa(\reg_file[23][18]~q ),
	.datab(\Mux13~7_combout ),
	.datac(\reg_file[31][18]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux13~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~8 .lut_mask = 16'hE2CC;
defparam \Mux13~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N28
cycloneive_lcell_comb \Mux13~0 (
// Equation(s):
// \Mux13~0_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[25][18]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & ((\reg_file[17][18]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[25][18]~q ),
	.datad(\reg_file[17][18]~q ),
	.cin(gnd),
	.combout(\Mux13~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~0 .lut_mask = 16'hB9A8;
defparam \Mux13~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N16
cycloneive_lcell_comb \Mux13~1 (
// Equation(s):
// \Mux13~1_combout  = (\prif.imemload_id [23] & ((\Mux13~0_combout  & ((\reg_file[29][18]~q ))) # (!\Mux13~0_combout  & (\reg_file[21][18]~q )))) # (!\prif.imemload_id [23] & (((\Mux13~0_combout ))))

	.dataa(\reg_file[21][18]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[29][18]~q ),
	.datad(\Mux13~0_combout ),
	.cin(gnd),
	.combout(\Mux13~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~1 .lut_mask = 16'hF388;
defparam \Mux13~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N14
cycloneive_lcell_comb \Mux13~2 (
// Equation(s):
// \Mux13~2_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[22][18]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[18][18]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[18][18]~q ),
	.datad(\reg_file[22][18]~q ),
	.cin(gnd),
	.combout(\Mux13~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~2 .lut_mask = 16'hBA98;
defparam \Mux13~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N24
cycloneive_lcell_comb \Mux13~3 (
// Equation(s):
// \Mux13~3_combout  = (\prif.imemload_id [24] & ((\Mux13~2_combout  & (\reg_file[30][18]~q )) # (!\Mux13~2_combout  & ((\reg_file[26][18]~q ))))) # (!\prif.imemload_id [24] & (((\Mux13~2_combout ))))

	.dataa(\reg_file[30][18]~q ),
	.datab(prifimemload_id_24),
	.datac(\Mux13~2_combout ),
	.datad(\reg_file[26][18]~q ),
	.cin(gnd),
	.combout(\Mux13~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~3 .lut_mask = 16'hBCB0;
defparam \Mux13~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N22
cycloneive_lcell_comb \reg_file[24][18]~feeder (
// Equation(s):
// \reg_file[24][18]~feeder_combout  = \reg_file_nxt[31][18]~83_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][18]~83_combout ),
	.cin(gnd),
	.combout(\reg_file[24][18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][18]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[24][18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N23
dffeas \reg_file[24][18] (
	.clk(!CLK),
	.d(\reg_file[24][18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][18] .is_wysiwyg = "true";
defparam \reg_file[24][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N2
cycloneive_lcell_comb \Mux13~5 (
// Equation(s):
// \Mux13~5_combout  = (\Mux13~4_combout  & (((\reg_file[28][18]~q ) # (!\prif.imemload_id [24])))) # (!\Mux13~4_combout  & (\reg_file[24][18]~q  & ((\prif.imemload_id [24]))))

	.dataa(\Mux13~4_combout ),
	.datab(\reg_file[24][18]~q ),
	.datac(\reg_file[28][18]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux13~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~5 .lut_mask = 16'hE4AA;
defparam \Mux13~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N22
cycloneive_lcell_comb \Mux13~6 (
// Equation(s):
// \Mux13~6_combout  = (\prif.imemload_id [22] & ((\Mux13~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\Mux13~5_combout  & !\prif.imemload_id [21]))))

	.dataa(\Mux13~3_combout ),
	.datab(prifimemload_id_22),
	.datac(\Mux13~5_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux13~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~6 .lut_mask = 16'hCCB8;
defparam \Mux13~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y27_N15
dffeas \reg_file[4][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][18] .is_wysiwyg = "true";
defparam \reg_file[4][18] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y27_N29
dffeas \reg_file[5][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][18] .is_wysiwyg = "true";
defparam \reg_file[5][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N28
cycloneive_lcell_comb \Mux13~10 (
// Equation(s):
// \Mux13~10_combout  = (\prif.imemload_id [21] & (((\reg_file[5][18]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[4][18]~q  & ((!\prif.imemload_id [22]))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[4][18]~q ),
	.datac(\reg_file[5][18]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux13~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~10 .lut_mask = 16'hAAE4;
defparam \Mux13~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N20
cycloneive_lcell_comb \Mux13~11 (
// Equation(s):
// \Mux13~11_combout  = (\prif.imemload_id [22] & ((\Mux13~10_combout  & (\reg_file[7][18]~q )) # (!\Mux13~10_combout  & ((\reg_file[6][18]~q ))))) # (!\prif.imemload_id [22] & (((\Mux13~10_combout ))))

	.dataa(\reg_file[7][18]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[6][18]~q ),
	.datad(\Mux13~10_combout ),
	.cin(gnd),
	.combout(\Mux13~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~11 .lut_mask = 16'hBBC0;
defparam \Mux13~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N31
dffeas \reg_file[12][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][18] .is_wysiwyg = "true";
defparam \reg_file[12][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N30
cycloneive_lcell_comb \Mux13~17 (
// Equation(s):
// \Mux13~17_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[13][18]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[12][18]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[12][18]~q ),
	.datad(\reg_file[13][18]~q ),
	.cin(gnd),
	.combout(\Mux13~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~17 .lut_mask = 16'hBA98;
defparam \Mux13~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N16
cycloneive_lcell_comb \Mux13~18 (
// Equation(s):
// \Mux13~18_combout  = (\prif.imemload_id [22] & ((\Mux13~17_combout  & (\reg_file[15][18]~q )) # (!\Mux13~17_combout  & ((\reg_file[14][18]~q ))))) # (!\prif.imemload_id [22] & (((\Mux13~17_combout ))))

	.dataa(\reg_file[15][18]~q ),
	.datab(\reg_file[14][18]~q ),
	.datac(prifimemload_id_22),
	.datad(\Mux13~17_combout ),
	.cin(gnd),
	.combout(\Mux13~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~18 .lut_mask = 16'hAFC0;
defparam \Mux13~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N31
dffeas \reg_file[3][18] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][18]~83_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][18]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][18] .is_wysiwyg = "true";
defparam \reg_file[3][18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N30
cycloneive_lcell_comb \Mux13~14 (
// Equation(s):
// \Mux13~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][18]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][18]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][18]~q ),
	.datad(\reg_file[1][18]~q ),
	.cin(gnd),
	.combout(\Mux13~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~14 .lut_mask = 16'hA280;
defparam \Mux13~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N14
cycloneive_lcell_comb \Mux13~15 (
// Equation(s):
// \Mux13~15_combout  = (\Mux13~14_combout ) # ((\reg_file[2][18]~q  & (\prif.imemload_id [22] & !\prif.imemload_id [21])))

	.dataa(\reg_file[2][18]~q ),
	.datab(prifimemload_id_22),
	.datac(\Mux13~14_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux13~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~15 .lut_mask = 16'hF0F8;
defparam \Mux13~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N12
cycloneive_lcell_comb \Mux13~13 (
// Equation(s):
// \Mux13~13_combout  = (\Mux13~12_combout  & ((\reg_file[11][18]~q ) # ((!\prif.imemload_id [21])))) # (!\Mux13~12_combout  & (((\reg_file[9][18]~q  & \prif.imemload_id [21]))))

	.dataa(\Mux13~12_combout ),
	.datab(\reg_file[11][18]~q ),
	.datac(\reg_file[9][18]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux13~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~13 .lut_mask = 16'hD8AA;
defparam \Mux13~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N24
cycloneive_lcell_comb \Mux13~16 (
// Equation(s):
// \Mux13~16_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\Mux13~13_combout ))) # (!\prif.imemload_id [24] & (\Mux13~15_combout ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux13~15_combout ),
	.datad(\Mux13~13_combout ),
	.cin(gnd),
	.combout(\Mux13~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux13~16 .lut_mask = 16'hDC98;
defparam \Mux13~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N26
cycloneive_lcell_comb \Mux14~0 (
// Equation(s):
// \Mux14~0_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24]) # (\reg_file[21][17]~q )))) # (!\prif.imemload_id [23] & (\reg_file[17][17]~q  & (!\prif.imemload_id [24])))

	.dataa(\reg_file[17][17]~q ),
	.datab(prifimemload_id_23),
	.datac(prifimemload_id_24),
	.datad(\reg_file[21][17]~q ),
	.cin(gnd),
	.combout(\Mux14~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~0 .lut_mask = 16'hCEC2;
defparam \Mux14~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N10
cycloneive_lcell_comb \Mux14~1 (
// Equation(s):
// \Mux14~1_combout  = (\Mux14~0_combout  & (((\reg_file[29][17]~q )) # (!\prif.imemload_id [24]))) # (!\Mux14~0_combout  & (\prif.imemload_id [24] & ((\reg_file[25][17]~q ))))

	.dataa(\Mux14~0_combout ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[29][17]~q ),
	.datad(\reg_file[25][17]~q ),
	.cin(gnd),
	.combout(\Mux14~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~1 .lut_mask = 16'hE6A2;
defparam \Mux14~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N6
cycloneive_lcell_comb \reg_file[26][17]~feeder (
// Equation(s):
// \reg_file[26][17]~feeder_combout  = \reg_file_nxt[31][17]~87_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][17]~87_combout ),
	.cin(gnd),
	.combout(\reg_file[26][17]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[26][17]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[26][17]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N7
dffeas \reg_file[26][17] (
	.clk(!CLK),
	.d(\reg_file[26][17]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][17] .is_wysiwyg = "true";
defparam \reg_file[26][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N6
cycloneive_lcell_comb \Mux14~2 (
// Equation(s):
// \Mux14~2_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[26][17]~q ))) # (!\prif.imemload_id [24] & (\reg_file[18][17]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[18][17]~q ),
	.datad(\reg_file[26][17]~q ),
	.cin(gnd),
	.combout(\Mux14~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~2 .lut_mask = 16'hDC98;
defparam \Mux14~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N26
cycloneive_lcell_comb \Mux14~3 (
// Equation(s):
// \Mux14~3_combout  = (\prif.imemload_id [23] & ((\Mux14~2_combout  & (\reg_file[30][17]~q )) # (!\Mux14~2_combout  & ((\reg_file[22][17]~q ))))) # (!\prif.imemload_id [23] & (((\Mux14~2_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[30][17]~q ),
	.datac(\reg_file[22][17]~q ),
	.datad(\Mux14~2_combout ),
	.cin(gnd),
	.combout(\Mux14~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~3 .lut_mask = 16'hDDA0;
defparam \Mux14~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N7
dffeas \reg_file[16][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][17] .is_wysiwyg = "true";
defparam \reg_file[16][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N16
cycloneive_lcell_comb \Mux14~4 (
// Equation(s):
// \Mux14~4_combout  = (\prif.imemload_id [24] & (((\reg_file[24][17]~q ) # (\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (\reg_file[16][17]~q  & ((!\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[16][17]~q ),
	.datac(\reg_file[24][17]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux14~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~4 .lut_mask = 16'hAAE4;
defparam \Mux14~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N26
cycloneive_lcell_comb \Mux14~5 (
// Equation(s):
// \Mux14~5_combout  = (\prif.imemload_id [23] & ((\Mux14~4_combout  & ((\reg_file[28][17]~q ))) # (!\Mux14~4_combout  & (\reg_file[20][17]~q )))) # (!\prif.imemload_id [23] & (((\Mux14~4_combout ))))

	.dataa(\reg_file[20][17]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[28][17]~q ),
	.datad(\Mux14~4_combout ),
	.cin(gnd),
	.combout(\Mux14~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~5 .lut_mask = 16'hF388;
defparam \Mux14~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N20
cycloneive_lcell_comb \Mux14~6 (
// Equation(s):
// \Mux14~6_combout  = (\prif.imemload_id [22] & ((\Mux14~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\Mux14~5_combout  & !\prif.imemload_id [21]))))

	.dataa(prifimemload_id_22),
	.datab(\Mux14~3_combout ),
	.datac(\Mux14~5_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux14~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~6 .lut_mask = 16'hAAD8;
defparam \Mux14~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N2
cycloneive_lcell_comb \Mux14~7 (
// Equation(s):
// \Mux14~7_combout  = (\prif.imemload_id [23] & ((\reg_file[23][17]~q ) # ((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (((\reg_file[19][17]~q  & !\prif.imemload_id [24]))))

	.dataa(\reg_file[23][17]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][17]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux14~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~7 .lut_mask = 16'hCCB8;
defparam \Mux14~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y34_N26
cycloneive_lcell_comb \Mux14~8 (
// Equation(s):
// \Mux14~8_combout  = (\Mux14~7_combout  & ((\reg_file[31][17]~q ) # ((!\prif.imemload_id [24])))) # (!\Mux14~7_combout  & (((\prif.imemload_id [24] & \reg_file[27][17]~q ))))

	.dataa(\Mux14~7_combout ),
	.datab(\reg_file[31][17]~q ),
	.datac(prifimemload_id_24),
	.datad(\reg_file[27][17]~q ),
	.cin(gnd),
	.combout(\Mux14~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~8 .lut_mask = 16'hDA8A;
defparam \Mux14~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N6
cycloneive_lcell_comb \Mux14~17 (
// Equation(s):
// \Mux14~17_combout  = (\prif.imemload_id [21] & ((\reg_file[13][17]~q ) # ((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (((\reg_file[12][17]~q  & !\prif.imemload_id [22]))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[13][17]~q ),
	.datac(\reg_file[12][17]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux14~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~17 .lut_mask = 16'hAAD8;
defparam \Mux14~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N18
cycloneive_lcell_comb \Mux14~18 (
// Equation(s):
// \Mux14~18_combout  = (\prif.imemload_id [22] & ((\Mux14~17_combout  & (\reg_file[15][17]~q )) # (!\Mux14~17_combout  & ((\reg_file[14][17]~q ))))) # (!\prif.imemload_id [22] & (((\Mux14~17_combout ))))

	.dataa(\reg_file[15][17]~q ),
	.datab(\reg_file[14][17]~q ),
	.datac(prifimemload_id_22),
	.datad(\Mux14~17_combout ),
	.cin(gnd),
	.combout(\Mux14~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~18 .lut_mask = 16'hAFC0;
defparam \Mux14~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N23
dffeas \reg_file[2][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~48_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[2][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[2][17] .is_wysiwyg = "true";
defparam \reg_file[2][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N22
cycloneive_lcell_comb \Mux14~15 (
// Equation(s):
// \Mux14~15_combout  = (\Mux14~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][17]~q  & !\prif.imemload_id [21])))

	.dataa(\Mux14~14_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][17]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux14~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~15 .lut_mask = 16'hAAEA;
defparam \Mux14~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N22
cycloneive_lcell_comb \Mux14~13 (
// Equation(s):
// \Mux14~13_combout  = (\Mux14~12_combout  & (((\reg_file[7][17]~q )) # (!\prif.imemload_id [22]))) # (!\Mux14~12_combout  & (\prif.imemload_id [22] & ((\reg_file[6][17]~q ))))

	.dataa(\Mux14~12_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[7][17]~q ),
	.datad(\reg_file[6][17]~q ),
	.cin(gnd),
	.combout(\Mux14~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~13 .lut_mask = 16'hE6A2;
defparam \Mux14~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N8
cycloneive_lcell_comb \Mux14~16 (
// Equation(s):
// \Mux14~16_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\Mux14~13_combout )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\Mux14~15_combout )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux14~15_combout ),
	.datad(\Mux14~13_combout ),
	.cin(gnd),
	.combout(\Mux14~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~16 .lut_mask = 16'hBA98;
defparam \Mux14~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N20
cycloneive_lcell_comb \Mux14~10 (
// Equation(s):
// \Mux14~10_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[10][17]~q ))) # (!\prif.imemload_id [22] & (\reg_file[8][17]~q ))))

	.dataa(\reg_file[8][17]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[10][17]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux14~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~10 .lut_mask = 16'hFC22;
defparam \Mux14~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y33_N19
dffeas \reg_file[11][17] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][17]~87_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][17]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][17] .is_wysiwyg = "true";
defparam \reg_file[11][17] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y33_N18
cycloneive_lcell_comb \Mux14~11 (
// Equation(s):
// \Mux14~11_combout  = (\Mux14~10_combout  & (((\reg_file[11][17]~q ) # (!\prif.imemload_id [21])))) # (!\Mux14~10_combout  & (\reg_file[9][17]~q  & ((\prif.imemload_id [21]))))

	.dataa(\reg_file[9][17]~q ),
	.datab(\Mux14~10_combout ),
	.datac(\reg_file[11][17]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux14~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux14~11 .lut_mask = 16'hE2CC;
defparam \Mux14~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N8
cycloneive_lcell_comb \Mux11~0 (
// Equation(s):
// \Mux11~0_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][20]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][20]~q )))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[25][20]~q ),
	.datac(\reg_file[17][20]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux11~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~0 .lut_mask = 16'hEE50;
defparam \Mux11~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N20
cycloneive_lcell_comb \Mux11~1 (
// Equation(s):
// \Mux11~1_combout  = (\Mux11~0_combout  & (((\reg_file[29][20]~q ) # (!\prif.imemload_id [23])))) # (!\Mux11~0_combout  & (\reg_file[21][20]~q  & (\prif.imemload_id [23])))

	.dataa(\Mux11~0_combout ),
	.datab(\reg_file[21][20]~q ),
	.datac(prifimemload_id_23),
	.datad(\reg_file[29][20]~q ),
	.cin(gnd),
	.combout(\Mux11~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~1 .lut_mask = 16'hEA4A;
defparam \Mux11~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N10
cycloneive_lcell_comb \Mux11~7 (
// Equation(s):
// \Mux11~7_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[27][20]~q ))) # (!\prif.imemload_id [24] & (\reg_file[19][20]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[19][20]~q ),
	.datad(\reg_file[27][20]~q ),
	.cin(gnd),
	.combout(\Mux11~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~7 .lut_mask = 16'hDC98;
defparam \Mux11~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N26
cycloneive_lcell_comb \Mux11~8 (
// Equation(s):
// \Mux11~8_combout  = (\Mux11~7_combout  & ((\reg_file[31][20]~q ) # ((!\prif.imemload_id [23])))) # (!\Mux11~7_combout  & (((\prif.imemload_id [23] & \reg_file[23][20]~q ))))

	.dataa(\Mux11~7_combout ),
	.datab(\reg_file[31][20]~q ),
	.datac(prifimemload_id_23),
	.datad(\reg_file[23][20]~q ),
	.cin(gnd),
	.combout(\Mux11~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~8 .lut_mask = 16'hDA8A;
defparam \Mux11~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N5
dffeas \reg_file[26][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][20] .is_wysiwyg = "true";
defparam \reg_file[26][20] .power_up = "low";
// synopsys translate_on

// Location: FF_X65_Y31_N19
dffeas \reg_file[18][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][20] .is_wysiwyg = "true";
defparam \reg_file[18][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N18
cycloneive_lcell_comb \Mux11~2 (
// Equation(s):
// \Mux11~2_combout  = (\prif.imemload_id [23] & ((\reg_file[22][20]~q ) # ((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (((\reg_file[18][20]~q  & !\prif.imemload_id [24]))))

	.dataa(\reg_file[22][20]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[18][20]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux11~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~2 .lut_mask = 16'hCCB8;
defparam \Mux11~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N10
cycloneive_lcell_comb \Mux11~3 (
// Equation(s):
// \Mux11~3_combout  = (\prif.imemload_id [24] & ((\Mux11~2_combout  & ((\reg_file[30][20]~q ))) # (!\Mux11~2_combout  & (\reg_file[26][20]~q )))) # (!\prif.imemload_id [24] & (((\Mux11~2_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[26][20]~q ),
	.datac(\reg_file[30][20]~q ),
	.datad(\Mux11~2_combout ),
	.cin(gnd),
	.combout(\Mux11~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~3 .lut_mask = 16'hF588;
defparam \Mux11~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N28
cycloneive_lcell_comb \Mux11~4 (
// Equation(s):
// \Mux11~4_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\reg_file[20][20]~q )) # (!\prif.imemload_id [23] & ((\reg_file[16][20]~q )))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[20][20]~q ),
	.datad(\reg_file[16][20]~q ),
	.cin(gnd),
	.combout(\Mux11~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~4 .lut_mask = 16'hD9C8;
defparam \Mux11~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N14
cycloneive_lcell_comb \Mux11~5 (
// Equation(s):
// \Mux11~5_combout  = (\prif.imemload_id [24] & ((\Mux11~4_combout  & ((\reg_file[28][20]~q ))) # (!\Mux11~4_combout  & (\reg_file[24][20]~q )))) # (!\prif.imemload_id [24] & (((\Mux11~4_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[24][20]~q ),
	.datac(\reg_file[28][20]~q ),
	.datad(\Mux11~4_combout ),
	.cin(gnd),
	.combout(\Mux11~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~5 .lut_mask = 16'hF588;
defparam \Mux11~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N28
cycloneive_lcell_comb \Mux11~6 (
// Equation(s):
// \Mux11~6_combout  = (\prif.imemload_id [22] & ((\Mux11~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((!\prif.imemload_id [21] & \Mux11~5_combout ))))

	.dataa(\Mux11~3_combout ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux11~5_combout ),
	.cin(gnd),
	.combout(\Mux11~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~6 .lut_mask = 16'hCBC8;
defparam \Mux11~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y31_N23
dffeas \reg_file[12][20] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][20]~89_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][20] .is_wysiwyg = "true";
defparam \reg_file[12][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y31_N22
cycloneive_lcell_comb \Mux11~17 (
// Equation(s):
// \Mux11~17_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[13][20]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[12][20]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[12][20]~q ),
	.datad(\reg_file[13][20]~q ),
	.cin(gnd),
	.combout(\Mux11~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~17 .lut_mask = 16'hBA98;
defparam \Mux11~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N14
cycloneive_lcell_comb \Mux11~18 (
// Equation(s):
// \Mux11~18_combout  = (\Mux11~17_combout  & ((\reg_file[15][20]~q ) # ((!\prif.imemload_id [22])))) # (!\Mux11~17_combout  & (((\prif.imemload_id [22] & \reg_file[14][20]~q ))))

	.dataa(\reg_file[15][20]~q ),
	.datab(\Mux11~17_combout ),
	.datac(prifimemload_id_22),
	.datad(\reg_file[14][20]~q ),
	.cin(gnd),
	.combout(\Mux11~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~18 .lut_mask = 16'hBC8C;
defparam \Mux11~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N22
cycloneive_lcell_comb \reg_file[6][20]~feeder (
// Equation(s):
// \reg_file[6][20]~feeder_combout  = \reg_file_nxt[31][20]~89_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][20]~89_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[6][20]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[6][20]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[6][20]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y28_N23
dffeas \reg_file[6][20] (
	.clk(!CLK),
	.d(\reg_file[6][20]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~42_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[6][20]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[6][20] .is_wysiwyg = "true";
defparam \reg_file[6][20] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N6
cycloneive_lcell_comb \Mux11~10 (
// Equation(s):
// \Mux11~10_combout  = (\prif.imemload_id [21] & ((\reg_file[5][20]~q ) # ((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (((\reg_file[4][20]~q  & !\prif.imemload_id [22]))))

	.dataa(\reg_file[5][20]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[4][20]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux11~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~10 .lut_mask = 16'hCCB8;
defparam \Mux11~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N12
cycloneive_lcell_comb \Mux11~11 (
// Equation(s):
// \Mux11~11_combout  = (\prif.imemload_id [22] & ((\Mux11~10_combout  & ((\reg_file[7][20]~q ))) # (!\Mux11~10_combout  & (\reg_file[6][20]~q )))) # (!\prif.imemload_id [22] & (((\Mux11~10_combout ))))

	.dataa(\reg_file[6][20]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[7][20]~q ),
	.datad(\Mux11~10_combout ),
	.cin(gnd),
	.combout(\Mux11~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~11 .lut_mask = 16'hF388;
defparam \Mux11~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N30
cycloneive_lcell_comb \Mux11~13 (
// Equation(s):
// \Mux11~13_combout  = (\Mux11~12_combout  & (((\reg_file[11][20]~q ) # (!\prif.imemload_id [21])))) # (!\Mux11~12_combout  & (\reg_file[9][20]~q  & ((\prif.imemload_id [21]))))

	.dataa(\Mux11~12_combout ),
	.datab(\reg_file[9][20]~q ),
	.datac(\reg_file[11][20]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux11~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~13 .lut_mask = 16'hE4AA;
defparam \Mux11~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N16
cycloneive_lcell_comb \Mux11~15 (
// Equation(s):
// \Mux11~15_combout  = (\Mux11~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][20]~q  & !\prif.imemload_id [21])))

	.dataa(\Mux11~14_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][20]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux11~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~15 .lut_mask = 16'hAAEA;
defparam \Mux11~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N10
cycloneive_lcell_comb \Mux11~16 (
// Equation(s):
// \Mux11~16_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\Mux11~13_combout )) # (!\prif.imemload_id [24] & ((\Mux11~15_combout )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux11~13_combout ),
	.datad(\Mux11~15_combout ),
	.cin(gnd),
	.combout(\Mux11~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux11~16 .lut_mask = 16'hD9C8;
defparam \Mux11~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N6
cycloneive_lcell_comb \Mux12~0 (
// Equation(s):
// \Mux12~0_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[21][19]~q ))) # (!\prif.imemload_id [23] & (\reg_file[17][19]~q ))))

	.dataa(\reg_file[17][19]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[21][19]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux12~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~0 .lut_mask = 16'hFC22;
defparam \Mux12~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N16
cycloneive_lcell_comb \Mux12~1 (
// Equation(s):
// \Mux12~1_combout  = (\Mux12~0_combout  & (((\reg_file[29][19]~q )) # (!\prif.imemload_id [24]))) # (!\Mux12~0_combout  & (\prif.imemload_id [24] & (\reg_file[25][19]~q )))

	.dataa(\Mux12~0_combout ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[25][19]~q ),
	.datad(\reg_file[29][19]~q ),
	.cin(gnd),
	.combout(\Mux12~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~1 .lut_mask = 16'hEA62;
defparam \Mux12~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N4
cycloneive_lcell_comb \Mux12~3 (
// Equation(s):
// \Mux12~3_combout  = (\Mux12~2_combout  & (((\reg_file[30][19]~q ) # (!\prif.imemload_id [23])))) # (!\Mux12~2_combout  & (\reg_file[22][19]~q  & (\prif.imemload_id [23])))

	.dataa(\Mux12~2_combout ),
	.datab(\reg_file[22][19]~q ),
	.datac(prifimemload_id_23),
	.datad(\reg_file[30][19]~q ),
	.cin(gnd),
	.combout(\Mux12~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~3 .lut_mask = 16'hEA4A;
defparam \Mux12~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N1
dffeas \reg_file[24][19] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][19]~86_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][19] .is_wysiwyg = "true";
defparam \reg_file[24][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N0
cycloneive_lcell_comb \Mux12~4 (
// Equation(s):
// \Mux12~4_combout  = (\prif.imemload_id [24] & (((\reg_file[24][19]~q ) # (\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (\reg_file[16][19]~q  & ((!\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[16][19]~q ),
	.datac(\reg_file[24][19]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux12~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~4 .lut_mask = 16'hAAE4;
defparam \Mux12~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N10
cycloneive_lcell_comb \Mux12~5 (
// Equation(s):
// \Mux12~5_combout  = (\prif.imemload_id [23] & ((\Mux12~4_combout  & ((\reg_file[28][19]~q ))) # (!\Mux12~4_combout  & (\reg_file[20][19]~q )))) # (!\prif.imemload_id [23] & (((\Mux12~4_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[20][19]~q ),
	.datac(\reg_file[28][19]~q ),
	.datad(\Mux12~4_combout ),
	.cin(gnd),
	.combout(\Mux12~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~5 .lut_mask = 16'hF588;
defparam \Mux12~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N14
cycloneive_lcell_comb \Mux12~6 (
// Equation(s):
// \Mux12~6_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\Mux12~3_combout )) # (!\prif.imemload_id [22] & ((\Mux12~5_combout )))))

	.dataa(prifimemload_id_21),
	.datab(\Mux12~3_combout ),
	.datac(\Mux12~5_combout ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux12~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~6 .lut_mask = 16'hEE50;
defparam \Mux12~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N14
cycloneive_lcell_comb \Mux12~7 (
// Equation(s):
// \Mux12~7_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\reg_file[23][19]~q )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\reg_file[19][19]~q )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[19][19]~q ),
	.datad(\reg_file[23][19]~q ),
	.cin(gnd),
	.combout(\Mux12~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~7 .lut_mask = 16'hBA98;
defparam \Mux12~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N0
cycloneive_lcell_comb \Mux12~8 (
// Equation(s):
// \Mux12~8_combout  = (\Mux12~7_combout  & ((\reg_file[31][19]~q ) # ((!\prif.imemload_id [24])))) # (!\Mux12~7_combout  & (((\reg_file[27][19]~q  & \prif.imemload_id [24]))))

	.dataa(\reg_file[31][19]~q ),
	.datab(\reg_file[27][19]~q ),
	.datac(\Mux12~7_combout ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux12~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~8 .lut_mask = 16'hACF0;
defparam \Mux12~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N24
cycloneive_lcell_comb \reg_file[11][19]~feeder (
// Equation(s):
// \reg_file[11][19]~feeder_combout  = \reg_file_nxt[31][19]~86_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][19]~86_combout ),
	.cin(gnd),
	.combout(\reg_file[11][19]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[11][19]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[11][19]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y33_N25
dffeas \reg_file[11][19] (
	.clk(!CLK),
	.d(\reg_file[11][19]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~37_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[11][19]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[11][19] .is_wysiwyg = "true";
defparam \reg_file[11][19] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y33_N24
cycloneive_lcell_comb \Mux12~10 (
// Equation(s):
// \Mux12~10_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[10][19]~q ))) # (!\prif.imemload_id [22] & (\reg_file[8][19]~q ))))

	.dataa(\reg_file[8][19]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[10][19]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux12~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~10 .lut_mask = 16'hFC22;
defparam \Mux12~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y32_N4
cycloneive_lcell_comb \Mux12~11 (
// Equation(s):
// \Mux12~11_combout  = (\prif.imemload_id [21] & ((\Mux12~10_combout  & (\reg_file[11][19]~q )) # (!\Mux12~10_combout  & ((\reg_file[9][19]~q ))))) # (!\prif.imemload_id [21] & (((\Mux12~10_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[11][19]~q ),
	.datac(\reg_file[9][19]~q ),
	.datad(\Mux12~10_combout ),
	.cin(gnd),
	.combout(\Mux12~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~11 .lut_mask = 16'hDDA0;
defparam \Mux12~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N20
cycloneive_lcell_comb \Mux12~17 (
// Equation(s):
// \Mux12~17_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[13][19]~q )) # (!\prif.imemload_id [21] & ((\reg_file[12][19]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[13][19]~q ),
	.datad(\reg_file[12][19]~q ),
	.cin(gnd),
	.combout(\Mux12~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~17 .lut_mask = 16'hD9C8;
defparam \Mux12~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N18
cycloneive_lcell_comb \Mux12~18 (
// Equation(s):
// \Mux12~18_combout  = (\Mux12~17_combout  & ((\reg_file[15][19]~q ) # ((!\prif.imemload_id [22])))) # (!\Mux12~17_combout  & (((\reg_file[14][19]~q  & \prif.imemload_id [22]))))

	.dataa(\Mux12~17_combout ),
	.datab(\reg_file[15][19]~q ),
	.datac(\reg_file[14][19]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux12~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~18 .lut_mask = 16'hD8AA;
defparam \Mux12~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N0
cycloneive_lcell_comb \Mux12~12 (
// Equation(s):
// \Mux12~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][19]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & ((\reg_file[4][19]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[5][19]~q ),
	.datad(\reg_file[4][19]~q ),
	.cin(gnd),
	.combout(\Mux12~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~12 .lut_mask = 16'hB9A8;
defparam \Mux12~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N30
cycloneive_lcell_comb \Mux12~13 (
// Equation(s):
// \Mux12~13_combout  = (\prif.imemload_id [22] & ((\Mux12~12_combout  & (\reg_file[7][19]~q )) # (!\Mux12~12_combout  & ((\reg_file[6][19]~q ))))) # (!\prif.imemload_id [22] & (((\Mux12~12_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[7][19]~q ),
	.datac(\reg_file[6][19]~q ),
	.datad(\Mux12~12_combout ),
	.cin(gnd),
	.combout(\Mux12~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~13 .lut_mask = 16'hDDA0;
defparam \Mux12~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N2
cycloneive_lcell_comb \Mux12~14 (
// Equation(s):
// \Mux12~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][19]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][19]~q ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[1][19]~q ),
	.datac(\reg_file[3][19]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux12~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~14 .lut_mask = 16'hA088;
defparam \Mux12~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N12
cycloneive_lcell_comb \Mux12~15 (
// Equation(s):
// \Mux12~15_combout  = (\Mux12~14_combout ) # ((!\prif.imemload_id [21] & (\reg_file[2][19]~q  & \prif.imemload_id [22])))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[2][19]~q ),
	.datac(\Mux12~14_combout ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux12~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~15 .lut_mask = 16'hF4F0;
defparam \Mux12~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y33_N18
cycloneive_lcell_comb \Mux12~16 (
// Equation(s):
// \Mux12~16_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\Mux12~13_combout )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & ((\Mux12~15_combout ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux12~13_combout ),
	.datad(\Mux12~15_combout ),
	.cin(gnd),
	.combout(\Mux12~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux12~16 .lut_mask = 16'hB9A8;
defparam \Mux12~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N16
cycloneive_lcell_comb \Mux9~0 (
// Equation(s):
// \Mux9~0_combout  = (\prif.imemload_id [24] & ((\reg_file[25][22]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[17][22]~q  & !\prif.imemload_id [23]))))

	.dataa(\reg_file[25][22]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[17][22]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux9~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~0 .lut_mask = 16'hCCB8;
defparam \Mux9~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N28
cycloneive_lcell_comb \Mux9~1 (
// Equation(s):
// \Mux9~1_combout  = (\prif.imemload_id [23] & ((\Mux9~0_combout  & (\reg_file[29][22]~q )) # (!\Mux9~0_combout  & ((\reg_file[21][22]~q ))))) # (!\prif.imemload_id [23] & (((\Mux9~0_combout ))))

	.dataa(\reg_file[29][22]~q ),
	.datab(\reg_file[21][22]~q ),
	.datac(prifimemload_id_23),
	.datad(\Mux9~0_combout ),
	.cin(gnd),
	.combout(\Mux9~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~1 .lut_mask = 16'hAFC0;
defparam \Mux9~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N30
cycloneive_lcell_comb \Mux9~7 (
// Equation(s):
// \Mux9~7_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[27][22]~q )) # (!\prif.imemload_id [24] & ((\reg_file[19][22]~q )))))

	.dataa(\reg_file[27][22]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][22]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux9~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~7 .lut_mask = 16'hEE30;
defparam \Mux9~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N0
cycloneive_lcell_comb \Mux9~8 (
// Equation(s):
// \Mux9~8_combout  = (\prif.imemload_id [23] & ((\Mux9~7_combout  & ((\reg_file[31][22]~q ))) # (!\Mux9~7_combout  & (\reg_file[23][22]~q )))) # (!\prif.imemload_id [23] & (\Mux9~7_combout ))

	.dataa(prifimemload_id_23),
	.datab(\Mux9~7_combout ),
	.datac(\reg_file[23][22]~q ),
	.datad(\reg_file[31][22]~q ),
	.cin(gnd),
	.combout(\Mux9~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~8 .lut_mask = 16'hEC64;
defparam \Mux9~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N26
cycloneive_lcell_comb \Mux9~2 (
// Equation(s):
// \Mux9~2_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[22][22]~q ))) # (!\prif.imemload_id [23] & (\reg_file[18][22]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[18][22]~q ),
	.datad(\reg_file[22][22]~q ),
	.cin(gnd),
	.combout(\Mux9~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~2 .lut_mask = 16'hDC98;
defparam \Mux9~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y30_N14
cycloneive_lcell_comb \Mux9~3 (
// Equation(s):
// \Mux9~3_combout  = (\prif.imemload_id [24] & ((\Mux9~2_combout  & ((\reg_file[30][22]~q ))) # (!\Mux9~2_combout  & (\reg_file[26][22]~q )))) # (!\prif.imemload_id [24] & (((\Mux9~2_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[26][22]~q ),
	.datac(\Mux9~2_combout ),
	.datad(\reg_file[30][22]~q ),
	.cin(gnd),
	.combout(\Mux9~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~3 .lut_mask = 16'hF858;
defparam \Mux9~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N23
dffeas \reg_file[16][22] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][22]~94_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][22]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][22] .is_wysiwyg = "true";
defparam \reg_file[16][22] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N22
cycloneive_lcell_comb \Mux9~4 (
// Equation(s):
// \Mux9~4_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[20][22]~q ))) # (!\prif.imemload_id [23] & (\reg_file[16][22]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[16][22]~q ),
	.datad(\reg_file[20][22]~q ),
	.cin(gnd),
	.combout(\Mux9~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~4 .lut_mask = 16'hDC98;
defparam \Mux9~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N14
cycloneive_lcell_comb \Mux9~5 (
// Equation(s):
// \Mux9~5_combout  = (\prif.imemload_id [24] & ((\Mux9~4_combout  & ((\reg_file[28][22]~q ))) # (!\Mux9~4_combout  & (\reg_file[24][22]~q )))) # (!\prif.imemload_id [24] & (((\Mux9~4_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[24][22]~q ),
	.datac(\reg_file[28][22]~q ),
	.datad(\Mux9~4_combout ),
	.cin(gnd),
	.combout(\Mux9~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~5 .lut_mask = 16'hF588;
defparam \Mux9~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N26
cycloneive_lcell_comb \Mux9~6 (
// Equation(s):
// \Mux9~6_combout  = (\prif.imemload_id [22] & ((\Mux9~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((\Mux9~5_combout  & !\prif.imemload_id [21]))))

	.dataa(\Mux9~3_combout ),
	.datab(prifimemload_id_22),
	.datac(\Mux9~5_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux9~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~6 .lut_mask = 16'hCCB8;
defparam \Mux9~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N8
cycloneive_lcell_comb \Mux9~17 (
// Equation(s):
// \Mux9~17_combout  = (\prif.imemload_id [21] & (((\reg_file[13][22]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[12][22]~q  & ((!\prif.imemload_id [22]))))

	.dataa(\reg_file[12][22]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[13][22]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux9~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~17 .lut_mask = 16'hCCE2;
defparam \Mux9~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N4
cycloneive_lcell_comb \Mux9~18 (
// Equation(s):
// \Mux9~18_combout  = (\prif.imemload_id [22] & ((\Mux9~17_combout  & ((\reg_file[15][22]~q ))) # (!\Mux9~17_combout  & (\reg_file[14][22]~q )))) # (!\prif.imemload_id [22] & (((\Mux9~17_combout ))))

	.dataa(\reg_file[14][22]~q ),
	.datab(prifimemload_id_22),
	.datac(\Mux9~17_combout ),
	.datad(\reg_file[15][22]~q ),
	.cin(gnd),
	.combout(\Mux9~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~18 .lut_mask = 16'hF838;
defparam \Mux9~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N8
cycloneive_lcell_comb \Mux9~10 (
// Equation(s):
// \Mux9~10_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[5][22]~q ))) # (!\prif.imemload_id [21] & (\reg_file[4][22]~q ))))

	.dataa(\reg_file[4][22]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[5][22]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux9~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~10 .lut_mask = 16'hFC22;
defparam \Mux9~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y30_N16
cycloneive_lcell_comb \Mux9~11 (
// Equation(s):
// \Mux9~11_combout  = (\prif.imemload_id [22] & ((\Mux9~10_combout  & (\reg_file[7][22]~q )) # (!\Mux9~10_combout  & ((\reg_file[6][22]~q ))))) # (!\prif.imemload_id [22] & (((\Mux9~10_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[7][22]~q ),
	.datac(\reg_file[6][22]~q ),
	.datad(\Mux9~10_combout ),
	.cin(gnd),
	.combout(\Mux9~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~11 .lut_mask = 16'hDDA0;
defparam \Mux9~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N16
cycloneive_lcell_comb \Mux9~12 (
// Equation(s):
// \Mux9~12_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[10][22]~q )) # (!\prif.imemload_id [22] & ((\reg_file[8][22]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[10][22]~q ),
	.datad(\reg_file[8][22]~q ),
	.cin(gnd),
	.combout(\Mux9~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~12 .lut_mask = 16'hD9C8;
defparam \Mux9~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N18
cycloneive_lcell_comb \Mux9~13 (
// Equation(s):
// \Mux9~13_combout  = (\prif.imemload_id [21] & ((\Mux9~12_combout  & ((\reg_file[11][22]~q ))) # (!\Mux9~12_combout  & (\reg_file[9][22]~q )))) # (!\prif.imemload_id [21] & (((\Mux9~12_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[9][22]~q ),
	.datac(\reg_file[11][22]~q ),
	.datad(\Mux9~12_combout ),
	.cin(gnd),
	.combout(\Mux9~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~13 .lut_mask = 16'hF588;
defparam \Mux9~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N18
cycloneive_lcell_comb \Mux9~14 (
// Equation(s):
// \Mux9~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][22]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][22]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][22]~q ),
	.datad(\reg_file[1][22]~q ),
	.cin(gnd),
	.combout(\Mux9~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~14 .lut_mask = 16'hA280;
defparam \Mux9~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N28
cycloneive_lcell_comb \Mux9~15 (
// Equation(s):
// \Mux9~15_combout  = (\Mux9~14_combout ) # ((\reg_file[2][22]~q  & (\prif.imemload_id [22] & !\prif.imemload_id [21])))

	.dataa(\reg_file[2][22]~q ),
	.datab(prifimemload_id_22),
	.datac(\Mux9~14_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux9~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~15 .lut_mask = 16'hF0F8;
defparam \Mux9~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N6
cycloneive_lcell_comb \Mux9~16 (
// Equation(s):
// \Mux9~16_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\Mux9~13_combout )) # (!\prif.imemload_id [24] & ((\Mux9~15_combout )))))

	.dataa(prifimemload_id_23),
	.datab(\Mux9~13_combout ),
	.datac(prifimemload_id_24),
	.datad(\Mux9~15_combout ),
	.cin(gnd),
	.combout(\Mux9~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux9~16 .lut_mask = 16'hE5E0;
defparam \Mux9~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N5
dffeas \reg_file[24][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][21] .is_wysiwyg = "true";
defparam \reg_file[24][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N4
cycloneive_lcell_comb \Mux10~4 (
// Equation(s):
// \Mux10~4_combout  = (\prif.imemload_id [24] & (((\reg_file[24][21]~q ) # (\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (\reg_file[16][21]~q  & ((!\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[16][21]~q ),
	.datac(\reg_file[24][21]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux10~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~4 .lut_mask = 16'hAAE4;
defparam \Mux10~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N30
cycloneive_lcell_comb \Mux10~5 (
// Equation(s):
// \Mux10~5_combout  = (\Mux10~4_combout  & (((\reg_file[28][21]~q ) # (!\prif.imemload_id [23])))) # (!\Mux10~4_combout  & (\reg_file[20][21]~q  & ((\prif.imemload_id [23]))))

	.dataa(\reg_file[20][21]~q ),
	.datab(\Mux10~4_combout ),
	.datac(\reg_file[28][21]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux10~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~5 .lut_mask = 16'hE2CC;
defparam \Mux10~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N10
cycloneive_lcell_comb \Mux10~2 (
// Equation(s):
// \Mux10~2_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[26][21]~q ))) # (!\prif.imemload_id [24] & (\reg_file[18][21]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[18][21]~q ),
	.datad(\reg_file[26][21]~q ),
	.cin(gnd),
	.combout(\Mux10~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~2 .lut_mask = 16'hDC98;
defparam \Mux10~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N26
cycloneive_lcell_comb \Mux10~3 (
// Equation(s):
// \Mux10~3_combout  = (\Mux10~2_combout  & (((\reg_file[30][21]~q ) # (!\prif.imemload_id [23])))) # (!\Mux10~2_combout  & (\reg_file[22][21]~q  & ((\prif.imemload_id [23]))))

	.dataa(\reg_file[22][21]~q ),
	.datab(\Mux10~2_combout ),
	.datac(\reg_file[30][21]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux10~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~3 .lut_mask = 16'hE2CC;
defparam \Mux10~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y32_N30
cycloneive_lcell_comb \Mux10~6 (
// Equation(s):
// \Mux10~6_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\Mux10~3_combout ))) # (!\prif.imemload_id [22] & (\Mux10~5_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\Mux10~5_combout ),
	.datac(\Mux10~3_combout ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux10~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~6 .lut_mask = 16'hFA44;
defparam \Mux10~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y29_N27
dffeas \reg_file[19][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[19][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[19][21] .is_wysiwyg = "true";
defparam \reg_file[19][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N26
cycloneive_lcell_comb \Mux10~7 (
// Equation(s):
// \Mux10~7_combout  = (\prif.imemload_id [23] & ((\reg_file[23][21]~q ) # ((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (((\reg_file[19][21]~q  & !\prif.imemload_id [24]))))

	.dataa(\reg_file[23][21]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][21]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux10~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~7 .lut_mask = 16'hCCB8;
defparam \Mux10~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y29_N14
cycloneive_lcell_comb \Mux10~8 (
// Equation(s):
// \Mux10~8_combout  = (\Mux10~7_combout  & ((\reg_file[31][21]~q ) # ((!\prif.imemload_id [24])))) # (!\Mux10~7_combout  & (((\reg_file[27][21]~q  & \prif.imemload_id [24]))))

	.dataa(\Mux10~7_combout ),
	.datab(\reg_file[31][21]~q ),
	.datac(\reg_file[27][21]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux10~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~8 .lut_mask = 16'hD8AA;
defparam \Mux10~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N18
cycloneive_lcell_comb \Mux10~0 (
// Equation(s):
// \Mux10~0_combout  = (\prif.imemload_id [23] & (((\reg_file[21][21]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[17][21]~q  & ((!\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[17][21]~q ),
	.datac(\reg_file[21][21]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux10~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~0 .lut_mask = 16'hAAE4;
defparam \Mux10~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N26
cycloneive_lcell_comb \Mux10~1 (
// Equation(s):
// \Mux10~1_combout  = (\Mux10~0_combout  & ((\reg_file[29][21]~q ) # ((!\prif.imemload_id [24])))) # (!\Mux10~0_combout  & (((\prif.imemload_id [24] & \reg_file[25][21]~q ))))

	.dataa(\Mux10~0_combout ),
	.datab(\reg_file[29][21]~q ),
	.datac(prifimemload_id_24),
	.datad(\reg_file[25][21]~q ),
	.cin(gnd),
	.combout(\Mux10~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~1 .lut_mask = 16'hDA8A;
defparam \Mux10~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N12
cycloneive_lcell_comb \Mux10~10 (
// Equation(s):
// \Mux10~10_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[10][21]~q )) # (!\prif.imemload_id [22] & ((\reg_file[8][21]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[10][21]~q ),
	.datad(\reg_file[8][21]~q ),
	.cin(gnd),
	.combout(\Mux10~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~10 .lut_mask = 16'hD9C8;
defparam \Mux10~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y35_N31
dffeas \reg_file[9][21] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][21]~88_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][21]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][21] .is_wysiwyg = "true";
defparam \reg_file[9][21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N30
cycloneive_lcell_comb \Mux10~11 (
// Equation(s):
// \Mux10~11_combout  = (\prif.imemload_id [21] & ((\Mux10~10_combout  & ((\reg_file[11][21]~q ))) # (!\Mux10~10_combout  & (\reg_file[9][21]~q )))) # (!\prif.imemload_id [21] & (\Mux10~10_combout ))

	.dataa(prifimemload_id_21),
	.datab(\Mux10~10_combout ),
	.datac(\reg_file[9][21]~q ),
	.datad(\reg_file[11][21]~q ),
	.cin(gnd),
	.combout(\Mux10~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~11 .lut_mask = 16'hEC64;
defparam \Mux10~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N6
cycloneive_lcell_comb \Mux10~17 (
// Equation(s):
// \Mux10~17_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[13][21]~q ))) # (!\prif.imemload_id [21] & (\reg_file[12][21]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[12][21]~q ),
	.datad(\reg_file[13][21]~q ),
	.cin(gnd),
	.combout(\Mux10~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~17 .lut_mask = 16'hDC98;
defparam \Mux10~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y31_N10
cycloneive_lcell_comb \Mux10~18 (
// Equation(s):
// \Mux10~18_combout  = (\Mux10~17_combout  & ((\reg_file[15][21]~q ) # ((!\prif.imemload_id [22])))) # (!\Mux10~17_combout  & (((\reg_file[14][21]~q  & \prif.imemload_id [22]))))

	.dataa(\reg_file[15][21]~q ),
	.datab(\reg_file[14][21]~q ),
	.datac(\Mux10~17_combout ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux10~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~18 .lut_mask = 16'hACF0;
defparam \Mux10~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N24
cycloneive_lcell_comb \Mux10~12 (
// Equation(s):
// \Mux10~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][21]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & ((\reg_file[4][21]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[5][21]~q ),
	.datad(\reg_file[4][21]~q ),
	.cin(gnd),
	.combout(\Mux10~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~12 .lut_mask = 16'hB9A8;
defparam \Mux10~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N30
cycloneive_lcell_comb \Mux10~13 (
// Equation(s):
// \Mux10~13_combout  = (\prif.imemload_id [22] & ((\Mux10~12_combout  & ((\reg_file[7][21]~q ))) # (!\Mux10~12_combout  & (\reg_file[6][21]~q )))) # (!\prif.imemload_id [22] & (((\Mux10~12_combout ))))

	.dataa(\reg_file[6][21]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[7][21]~q ),
	.datad(\Mux10~12_combout ),
	.cin(gnd),
	.combout(\Mux10~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~13 .lut_mask = 16'hF388;
defparam \Mux10~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y33_N18
cycloneive_lcell_comb \Mux10~14 (
// Equation(s):
// \Mux10~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][21]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][21]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[1][21]~q ),
	.datad(\reg_file[3][21]~q ),
	.cin(gnd),
	.combout(\Mux10~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~14 .lut_mask = 16'hC840;
defparam \Mux10~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N0
cycloneive_lcell_comb \Mux10~15 (
// Equation(s):
// \Mux10~15_combout  = (\Mux10~14_combout ) # ((!\prif.imemload_id [21] & (\prif.imemload_id [22] & \reg_file[2][21]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][21]~q ),
	.datad(\Mux10~14_combout ),
	.cin(gnd),
	.combout(\Mux10~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~15 .lut_mask = 16'hFF40;
defparam \Mux10~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N26
cycloneive_lcell_comb \Mux10~16 (
// Equation(s):
// \Mux10~16_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\Mux10~13_combout )) # (!\prif.imemload_id [23] & ((\Mux10~15_combout )))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\Mux10~13_combout ),
	.datad(\Mux10~15_combout ),
	.cin(gnd),
	.combout(\Mux10~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux10~16 .lut_mask = 16'hD9C8;
defparam \Mux10~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N18
cycloneive_lcell_comb \Mux7~7 (
// Equation(s):
// \Mux7~7_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & ((\reg_file[27][24]~q ))) # (!\prif.imemload_id [24] & (\reg_file[19][24]~q ))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[19][24]~q ),
	.datad(\reg_file[27][24]~q ),
	.cin(gnd),
	.combout(\Mux7~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~7 .lut_mask = 16'hDC98;
defparam \Mux7~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y32_N2
cycloneive_lcell_comb \Mux7~8 (
// Equation(s):
// \Mux7~8_combout  = (\prif.imemload_id [23] & ((\Mux7~7_combout  & (\reg_file[31][24]~q )) # (!\Mux7~7_combout  & ((\reg_file[23][24]~q ))))) # (!\prif.imemload_id [23] & (((\Mux7~7_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[31][24]~q ),
	.datac(\Mux7~7_combout ),
	.datad(\reg_file[23][24]~q ),
	.cin(gnd),
	.combout(\Mux7~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~8 .lut_mask = 16'hDAD0;
defparam \Mux7~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y30_N8
cycloneive_lcell_comb \Mux7~0 (
// Equation(s):
// \Mux7~0_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[25][24]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & ((\reg_file[17][24]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[25][24]~q ),
	.datad(\reg_file[17][24]~q ),
	.cin(gnd),
	.combout(\Mux7~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~0 .lut_mask = 16'hB9A8;
defparam \Mux7~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N8
cycloneive_lcell_comb \Mux7~1 (
// Equation(s):
// \Mux7~1_combout  = (\prif.imemload_id [23] & ((\Mux7~0_combout  & (\reg_file[29][24]~q )) # (!\Mux7~0_combout  & ((\reg_file[21][24]~q ))))) # (!\prif.imemload_id [23] & (((\Mux7~0_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[29][24]~q ),
	.datac(\Mux7~0_combout ),
	.datad(\reg_file[21][24]~q ),
	.cin(gnd),
	.combout(\Mux7~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~1 .lut_mask = 16'hDAD0;
defparam \Mux7~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N14
cycloneive_lcell_comb \reg_file[30][24]~feeder (
// Equation(s):
// \reg_file[30][24]~feeder_combout  = \reg_file_nxt[31][24]~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][24]~84_combout ),
	.cin(gnd),
	.combout(\reg_file[30][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[30][24]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[30][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y32_N15
dffeas \reg_file[30][24] (
	.clk(!CLK),
	.d(\reg_file[30][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~25_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[30][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[30][24] .is_wysiwyg = "true";
defparam \reg_file[30][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N10
cycloneive_lcell_comb \Mux7~3 (
// Equation(s):
// \Mux7~3_combout  = (\Mux7~2_combout  & ((\reg_file[30][24]~q ) # ((!\prif.imemload_id [24])))) # (!\Mux7~2_combout  & (((\reg_file[26][24]~q  & \prif.imemload_id [24]))))

	.dataa(\Mux7~2_combout ),
	.datab(\reg_file[30][24]~q ),
	.datac(\reg_file[26][24]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux7~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~3 .lut_mask = 16'hD8AA;
defparam \Mux7~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N8
cycloneive_lcell_comb \reg_file[24][24]~feeder (
// Equation(s):
// \reg_file[24][24]~feeder_combout  = \reg_file_nxt[31][24]~84_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][24]~84_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[24][24]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[24][24]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[24][24]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y33_N9
dffeas \reg_file[24][24] (
	.clk(!CLK),
	.d(\reg_file[24][24]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][24]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][24] .is_wysiwyg = "true";
defparam \reg_file[24][24] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N6
cycloneive_lcell_comb \Mux7~5 (
// Equation(s):
// \Mux7~5_combout  = (\Mux7~4_combout  & (((\reg_file[28][24]~q ) # (!\prif.imemload_id [24])))) # (!\Mux7~4_combout  & (\reg_file[24][24]~q  & ((\prif.imemload_id [24]))))

	.dataa(\Mux7~4_combout ),
	.datab(\reg_file[24][24]~q ),
	.datac(\reg_file[28][24]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux7~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~5 .lut_mask = 16'hE4AA;
defparam \Mux7~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N16
cycloneive_lcell_comb \Mux7~6 (
// Equation(s):
// \Mux7~6_combout  = (\prif.imemload_id [22] & ((\prif.imemload_id [21]) # ((\Mux7~3_combout )))) # (!\prif.imemload_id [22] & (!\prif.imemload_id [21] & ((\Mux7~5_combout ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\Mux7~3_combout ),
	.datad(\Mux7~5_combout ),
	.cin(gnd),
	.combout(\Mux7~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~6 .lut_mask = 16'hB9A8;
defparam \Mux7~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N14
cycloneive_lcell_comb \Mux7~17 (
// Equation(s):
// \Mux7~17_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[13][24]~q ))) # (!\prif.imemload_id [21] & (\reg_file[12][24]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[12][24]~q ),
	.datad(\reg_file[13][24]~q ),
	.cin(gnd),
	.combout(\Mux7~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~17 .lut_mask = 16'hDC98;
defparam \Mux7~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X61_Y32_N22
cycloneive_lcell_comb \Mux7~18 (
// Equation(s):
// \Mux7~18_combout  = (\prif.imemload_id [22] & ((\Mux7~17_combout  & (\reg_file[15][24]~q )) # (!\Mux7~17_combout  & ((\reg_file[14][24]~q ))))) # (!\prif.imemload_id [22] & (((\Mux7~17_combout ))))

	.dataa(\reg_file[15][24]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[14][24]~q ),
	.datad(\Mux7~17_combout ),
	.cin(gnd),
	.combout(\Mux7~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~18 .lut_mask = 16'hBBC0;
defparam \Mux7~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y27_N16
cycloneive_lcell_comb \Mux7~10 (
// Equation(s):
// \Mux7~10_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][24]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & ((\reg_file[4][24]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[5][24]~q ),
	.datad(\reg_file[4][24]~q ),
	.cin(gnd),
	.combout(\Mux7~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~10 .lut_mask = 16'hB9A8;
defparam \Mux7~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N4
cycloneive_lcell_comb \Mux7~11 (
// Equation(s):
// \Mux7~11_combout  = (\prif.imemload_id [22] & ((\Mux7~10_combout  & (\reg_file[7][24]~q )) # (!\Mux7~10_combout  & ((\reg_file[6][24]~q ))))) # (!\prif.imemload_id [22] & (((\Mux7~10_combout ))))

	.dataa(\reg_file[7][24]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[6][24]~q ),
	.datad(\Mux7~10_combout ),
	.cin(gnd),
	.combout(\Mux7~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~11 .lut_mask = 16'hBBC0;
defparam \Mux7~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N10
cycloneive_lcell_comb \Mux7~13 (
// Equation(s):
// \Mux7~13_combout  = (\Mux7~12_combout  & (((\reg_file[11][24]~q ) # (!\prif.imemload_id [21])))) # (!\Mux7~12_combout  & (\reg_file[9][24]~q  & ((\prif.imemload_id [21]))))

	.dataa(\Mux7~12_combout ),
	.datab(\reg_file[9][24]~q ),
	.datac(\reg_file[11][24]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux7~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~13 .lut_mask = 16'hE4AA;
defparam \Mux7~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N28
cycloneive_lcell_comb \Mux7~15 (
// Equation(s):
// \Mux7~15_combout  = (\Mux7~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][24]~q  & !\prif.imemload_id [21])))

	.dataa(\Mux7~14_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[2][24]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux7~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~15 .lut_mask = 16'hAAEA;
defparam \Mux7~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N8
cycloneive_lcell_comb \Mux7~16 (
// Equation(s):
// \Mux7~16_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\Mux7~13_combout )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & ((\Mux7~15_combout ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\Mux7~13_combout ),
	.datad(\Mux7~15_combout ),
	.cin(gnd),
	.combout(\Mux7~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux7~16 .lut_mask = 16'hB9A8;
defparam \Mux7~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N30
cycloneive_lcell_comb \Mux8~2 (
// Equation(s):
// \Mux8~2_combout  = (\prif.imemload_id [24] & ((\reg_file[26][23]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[18][23]~q  & !\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[26][23]~q ),
	.datac(\reg_file[18][23]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux8~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~2 .lut_mask = 16'hAAD8;
defparam \Mux8~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N22
cycloneive_lcell_comb \Mux8~3 (
// Equation(s):
// \Mux8~3_combout  = (\Mux8~2_combout  & (((\reg_file[30][23]~q ) # (!\prif.imemload_id [23])))) # (!\Mux8~2_combout  & (\reg_file[22][23]~q  & (\prif.imemload_id [23])))

	.dataa(\reg_file[22][23]~q ),
	.datab(\Mux8~2_combout ),
	.datac(prifimemload_id_23),
	.datad(\reg_file[30][23]~q ),
	.cin(gnd),
	.combout(\Mux8~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~3 .lut_mask = 16'hEC2C;
defparam \Mux8~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N15
dffeas \reg_file[20][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][23] .is_wysiwyg = "true";
defparam \reg_file[20][23] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N17
dffeas \reg_file[16][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][23] .is_wysiwyg = "true";
defparam \reg_file[16][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N16
cycloneive_lcell_comb \Mux8~4 (
// Equation(s):
// \Mux8~4_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[24][23]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[16][23]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[16][23]~q ),
	.datad(\reg_file[24][23]~q ),
	.cin(gnd),
	.combout(\Mux8~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~4 .lut_mask = 16'hBA98;
defparam \Mux8~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N16
cycloneive_lcell_comb \Mux8~5 (
// Equation(s):
// \Mux8~5_combout  = (\prif.imemload_id [23] & ((\Mux8~4_combout  & ((\reg_file[28][23]~q ))) # (!\Mux8~4_combout  & (\reg_file[20][23]~q )))) # (!\prif.imemload_id [23] & (((\Mux8~4_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[20][23]~q ),
	.datac(\reg_file[28][23]~q ),
	.datad(\Mux8~4_combout ),
	.cin(gnd),
	.combout(\Mux8~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~5 .lut_mask = 16'hF588;
defparam \Mux8~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N24
cycloneive_lcell_comb \Mux8~6 (
// Equation(s):
// \Mux8~6_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\Mux8~3_combout )) # (!\prif.imemload_id [22] & ((\Mux8~5_combout )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux8~3_combout ),
	.datad(\Mux8~5_combout ),
	.cin(gnd),
	.combout(\Mux8~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~6 .lut_mask = 16'hD9C8;
defparam \Mux8~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N22
cycloneive_lcell_comb \reg_file[17][23]~feeder (
// Equation(s):
// \reg_file[17][23]~feeder_combout  = \reg_file_nxt[31][23]~82_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][23]~82_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[17][23]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[17][23]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[17][23]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y30_N23
dffeas \reg_file[17][23] (
	.clk(!CLK),
	.d(\reg_file[17][23]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~18_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[17][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[17][23] .is_wysiwyg = "true";
defparam \reg_file[17][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N12
cycloneive_lcell_comb \Mux8~0 (
// Equation(s):
// \Mux8~0_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\reg_file[21][23]~q )) # (!\prif.imemload_id [23] & ((\reg_file[17][23]~q )))))

	.dataa(\reg_file[21][23]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[17][23]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux8~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~0 .lut_mask = 16'hEE30;
defparam \Mux8~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N26
cycloneive_lcell_comb \Mux8~1 (
// Equation(s):
// \Mux8~1_combout  = (\Mux8~0_combout  & (((\reg_file[29][23]~q )) # (!\prif.imemload_id [24]))) # (!\Mux8~0_combout  & (\prif.imemload_id [24] & ((\reg_file[25][23]~q ))))

	.dataa(\Mux8~0_combout ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[29][23]~q ),
	.datad(\reg_file[25][23]~q ),
	.cin(gnd),
	.combout(\Mux8~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~1 .lut_mask = 16'hE6A2;
defparam \Mux8~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N6
cycloneive_lcell_comb \Mux8~7 (
// Equation(s):
// \Mux8~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][23]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][23]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][23]~q ),
	.datad(\reg_file[23][23]~q ),
	.cin(gnd),
	.combout(\Mux8~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~7 .lut_mask = 16'hDC98;
defparam \Mux8~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N22
cycloneive_lcell_comb \Mux8~8 (
// Equation(s):
// \Mux8~8_combout  = (\prif.imemload_id [24] & ((\Mux8~7_combout  & (\reg_file[31][23]~q )) # (!\Mux8~7_combout  & ((\reg_file[27][23]~q ))))) # (!\prif.imemload_id [24] & (((\Mux8~7_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[31][23]~q ),
	.datac(\reg_file[27][23]~q ),
	.datad(\Mux8~7_combout ),
	.cin(gnd),
	.combout(\Mux8~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~8 .lut_mask = 16'hDDA0;
defparam \Mux8~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N24
cycloneive_lcell_comb \Mux8~14 (
// Equation(s):
// \Mux8~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][23]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][23]~q ))))

	.dataa(\reg_file[1][23]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][23]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux8~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~14 .lut_mask = 16'hE200;
defparam \Mux8~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N2
cycloneive_lcell_comb \Mux8~15 (
// Equation(s):
// \Mux8~15_combout  = (\Mux8~14_combout ) # ((\reg_file[2][23]~q  & (\prif.imemload_id [22] & !\prif.imemload_id [21])))

	.dataa(\reg_file[2][23]~q ),
	.datab(prifimemload_id_22),
	.datac(\Mux8~14_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux8~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~15 .lut_mask = 16'hF0F8;
defparam \Mux8~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N16
cycloneive_lcell_comb \Mux8~12 (
// Equation(s):
// \Mux8~12_combout  = (\prif.imemload_id [21] & ((\reg_file[5][23]~q ) # ((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (((\reg_file[4][23]~q  & !\prif.imemload_id [22]))))

	.dataa(\reg_file[5][23]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[4][23]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux8~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~12 .lut_mask = 16'hCCB8;
defparam \Mux8~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N12
cycloneive_lcell_comb \Mux8~13 (
// Equation(s):
// \Mux8~13_combout  = (\Mux8~12_combout  & (((\reg_file[7][23]~q ) # (!\prif.imemload_id [22])))) # (!\Mux8~12_combout  & (\reg_file[6][23]~q  & ((\prif.imemload_id [22]))))

	.dataa(\reg_file[6][23]~q ),
	.datab(\reg_file[7][23]~q ),
	.datac(\Mux8~12_combout ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux8~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~13 .lut_mask = 16'hCAF0;
defparam \Mux8~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N20
cycloneive_lcell_comb \Mux8~16 (
// Equation(s):
// \Mux8~16_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\Mux8~13_combout ))) # (!\prif.imemload_id [23] & (\Mux8~15_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\Mux8~15_combout ),
	.datac(prifimemload_id_23),
	.datad(\Mux8~13_combout ),
	.cin(gnd),
	.combout(\Mux8~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~16 .lut_mask = 16'hF4A4;
defparam \Mux8~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N1
dffeas \reg_file[9][23] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][23]~82_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][23]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][23] .is_wysiwyg = "true";
defparam \reg_file[9][23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N20
cycloneive_lcell_comb \Mux8~10 (
// Equation(s):
// \Mux8~10_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[10][23]~q ))) # (!\prif.imemload_id [22] & (\reg_file[8][23]~q ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[8][23]~q ),
	.datac(\reg_file[10][23]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux8~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~10 .lut_mask = 16'hFA44;
defparam \Mux8~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N0
cycloneive_lcell_comb \Mux8~11 (
// Equation(s):
// \Mux8~11_combout  = (\prif.imemload_id [21] & ((\Mux8~10_combout  & (\reg_file[11][23]~q )) # (!\Mux8~10_combout  & ((\reg_file[9][23]~q ))))) # (!\prif.imemload_id [21] & (((\Mux8~10_combout ))))

	.dataa(\reg_file[11][23]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[9][23]~q ),
	.datad(\Mux8~10_combout ),
	.cin(gnd),
	.combout(\Mux8~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~11 .lut_mask = 16'hBBC0;
defparam \Mux8~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N0
cycloneive_lcell_comb \Mux8~17 (
// Equation(s):
// \Mux8~17_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[13][23]~q )) # (!\prif.imemload_id [21] & ((\reg_file[12][23]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[13][23]~q ),
	.datad(\reg_file[12][23]~q ),
	.cin(gnd),
	.combout(\Mux8~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~17 .lut_mask = 16'hD9C8;
defparam \Mux8~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N26
cycloneive_lcell_comb \Mux8~18 (
// Equation(s):
// \Mux8~18_combout  = (\prif.imemload_id [22] & ((\Mux8~17_combout  & (\reg_file[15][23]~q )) # (!\Mux8~17_combout  & ((\reg_file[14][23]~q ))))) # (!\prif.imemload_id [22] & (((\Mux8~17_combout ))))

	.dataa(\reg_file[15][23]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[14][23]~q ),
	.datad(\Mux8~17_combout ),
	.cin(gnd),
	.combout(\Mux8~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux8~18 .lut_mask = 16'hBBC0;
defparam \Mux8~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N20
cycloneive_lcell_comb \Mux0~0 (
// Equation(s):
// \Mux0~0_combout  = (\prif.imemload_id [23] & (((\reg_file[21][31]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[17][31]~q  & ((!\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[17][31]~q ),
	.datac(\reg_file[21][31]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~0 .lut_mask = 16'hAAE4;
defparam \Mux0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N28
cycloneive_lcell_comb \Mux0~1 (
// Equation(s):
// \Mux0~1_combout  = (\prif.imemload_id [24] & ((\Mux0~0_combout  & ((\reg_file[29][31]~q ))) # (!\Mux0~0_combout  & (\reg_file[25][31]~q )))) # (!\prif.imemload_id [24] & (((\Mux0~0_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[25][31]~q ),
	.datac(\reg_file[29][31]~q ),
	.datad(\Mux0~0_combout ),
	.cin(gnd),
	.combout(\Mux0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~1 .lut_mask = 16'hF588;
defparam \Mux0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y26_N8
cycloneive_lcell_comb \Mux0~7 (
// Equation(s):
// \Mux0~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][31]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][31]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][31]~q ),
	.datad(\reg_file[23][31]~q ),
	.cin(gnd),
	.combout(\Mux0~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~7 .lut_mask = 16'hDC98;
defparam \Mux0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N22
cycloneive_lcell_comb \Mux0~8 (
// Equation(s):
// \Mux0~8_combout  = (\Mux0~7_combout  & (((\reg_file[31][31]~q )) # (!\prif.imemload_id [24]))) # (!\Mux0~7_combout  & (\prif.imemload_id [24] & ((\reg_file[27][31]~q ))))

	.dataa(\Mux0~7_combout ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[31][31]~q ),
	.datad(\reg_file[27][31]~q ),
	.cin(gnd),
	.combout(\Mux0~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~8 .lut_mask = 16'hE6A2;
defparam \Mux0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N21
dffeas \reg_file[22][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][31] .is_wysiwyg = "true";
defparam \reg_file[22][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N20
cycloneive_lcell_comb \Mux0~3 (
// Equation(s):
// \Mux0~3_combout  = (\Mux0~2_combout  & (((\reg_file[30][31]~q )) # (!\prif.imemload_id [23]))) # (!\Mux0~2_combout  & (\prif.imemload_id [23] & (\reg_file[22][31]~q )))

	.dataa(\Mux0~2_combout ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[22][31]~q ),
	.datad(\reg_file[30][31]~q ),
	.cin(gnd),
	.combout(\Mux0~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~3 .lut_mask = 16'hEA62;
defparam \Mux0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y33_N1
dffeas \reg_file[20][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][31] .is_wysiwyg = "true";
defparam \reg_file[20][31] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N7
dffeas \reg_file[16][31] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][31]~69_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][31]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][31] .is_wysiwyg = "true";
defparam \reg_file[16][31] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N6
cycloneive_lcell_comb \Mux0~4 (
// Equation(s):
// \Mux0~4_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[24][31]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[16][31]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[16][31]~q ),
	.datad(\reg_file[24][31]~q ),
	.cin(gnd),
	.combout(\Mux0~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~4 .lut_mask = 16'hBA98;
defparam \Mux0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N22
cycloneive_lcell_comb \Mux0~5 (
// Equation(s):
// \Mux0~5_combout  = (\prif.imemload_id [23] & ((\Mux0~4_combout  & ((\reg_file[28][31]~q ))) # (!\Mux0~4_combout  & (\reg_file[20][31]~q )))) # (!\prif.imemload_id [23] & (((\Mux0~4_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[20][31]~q ),
	.datac(\Mux0~4_combout ),
	.datad(\reg_file[28][31]~q ),
	.cin(gnd),
	.combout(\Mux0~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~5 .lut_mask = 16'hF858;
defparam \Mux0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y34_N10
cycloneive_lcell_comb \Mux0~6 (
// Equation(s):
// \Mux0~6_combout  = (\prif.imemload_id [22] & ((\prif.imemload_id [21]) # ((\Mux0~3_combout )))) # (!\prif.imemload_id [22] & (!\prif.imemload_id [21] & ((\Mux0~5_combout ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\Mux0~3_combout ),
	.datad(\Mux0~5_combout ),
	.cin(gnd),
	.combout(\Mux0~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~6 .lut_mask = 16'hB9A8;
defparam \Mux0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N24
cycloneive_lcell_comb \Mux0~17 (
// Equation(s):
// \Mux0~17_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[13][31]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & ((\reg_file[12][31]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[13][31]~q ),
	.datad(\reg_file[12][31]~q ),
	.cin(gnd),
	.combout(\Mux0~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~17 .lut_mask = 16'hB9A8;
defparam \Mux0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y26_N24
cycloneive_lcell_comb \Mux0~18 (
// Equation(s):
// \Mux0~18_combout  = (\prif.imemload_id [22] & ((\Mux0~17_combout  & (\reg_file[15][31]~q )) # (!\Mux0~17_combout  & ((\reg_file[14][31]~q ))))) # (!\prif.imemload_id [22] & (((\Mux0~17_combout ))))

	.dataa(\reg_file[15][31]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[14][31]~q ),
	.datad(\Mux0~17_combout ),
	.cin(gnd),
	.combout(\Mux0~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~18 .lut_mask = 16'hBBC0;
defparam \Mux0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N0
cycloneive_lcell_comb \Mux0~10 (
// Equation(s):
// \Mux0~10_combout  = (\prif.imemload_id [22] & (((\reg_file[10][31]~q ) # (\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (\reg_file[8][31]~q  & ((!\prif.imemload_id [21]))))

	.dataa(\reg_file[8][31]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[10][31]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux0~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~10 .lut_mask = 16'hCCE2;
defparam \Mux0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N12
cycloneive_lcell_comb \Mux0~11 (
// Equation(s):
// \Mux0~11_combout  = (\Mux0~10_combout  & ((\reg_file[11][31]~q ) # ((!\prif.imemload_id [21])))) # (!\Mux0~10_combout  & (((\reg_file[9][31]~q  & \prif.imemload_id [21]))))

	.dataa(\reg_file[11][31]~q ),
	.datab(\Mux0~10_combout ),
	.datac(\reg_file[9][31]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux0~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~11 .lut_mask = 16'hB8CC;
defparam \Mux0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N22
cycloneive_lcell_comb \Mux0~12 (
// Equation(s):
// \Mux0~12_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[5][31]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[4][31]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[4][31]~q ),
	.datad(\reg_file[5][31]~q ),
	.cin(gnd),
	.combout(\Mux0~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~12 .lut_mask = 16'hBA98;
defparam \Mux0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N14
cycloneive_lcell_comb \Mux0~13 (
// Equation(s):
// \Mux0~13_combout  = (\prif.imemload_id [22] & ((\Mux0~12_combout  & ((\reg_file[7][31]~q ))) # (!\Mux0~12_combout  & (\reg_file[6][31]~q )))) # (!\prif.imemload_id [22] & (((\Mux0~12_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[6][31]~q ),
	.datac(\reg_file[7][31]~q ),
	.datad(\Mux0~12_combout ),
	.cin(gnd),
	.combout(\Mux0~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~13 .lut_mask = 16'hF588;
defparam \Mux0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N20
cycloneive_lcell_comb \Mux0~14 (
// Equation(s):
// \Mux0~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][31]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][31]~q ))))

	.dataa(\reg_file[1][31]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][31]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux0~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~14 .lut_mask = 16'hE200;
defparam \Mux0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N0
cycloneive_lcell_comb \Mux0~15 (
// Equation(s):
// \Mux0~15_combout  = (\Mux0~14_combout ) # ((\prif.imemload_id [22] & (!\prif.imemload_id [21] & \reg_file[2][31]~q )))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\Mux0~14_combout ),
	.datad(\reg_file[2][31]~q ),
	.cin(gnd),
	.combout(\Mux0~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~15 .lut_mask = 16'hF2F0;
defparam \Mux0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y34_N2
cycloneive_lcell_comb \Mux0~16 (
// Equation(s):
// \Mux0~16_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\Mux0~13_combout )) # (!\prif.imemload_id [23] & ((\Mux0~15_combout )))))

	.dataa(prifimemload_id_24),
	.datab(\Mux0~13_combout ),
	.datac(prifimemload_id_23),
	.datad(\Mux0~15_combout ),
	.cin(gnd),
	.combout(\Mux0~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux0~16 .lut_mask = 16'hE5E0;
defparam \Mux0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N8
cycloneive_lcell_comb \Mux1~0 (
// Equation(s):
// \Mux1~0_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][30]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][30]~q )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[25][30]~q ),
	.datad(\reg_file[17][30]~q ),
	.cin(gnd),
	.combout(\Mux1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~0 .lut_mask = 16'hD9C8;
defparam \Mux1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N8
cycloneive_lcell_comb \Mux1~1 (
// Equation(s):
// \Mux1~1_combout  = (\prif.imemload_id [23] & ((\Mux1~0_combout  & ((\reg_file[29][30]~q ))) # (!\Mux1~0_combout  & (\reg_file[21][30]~q )))) # (!\prif.imemload_id [23] & (((\Mux1~0_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[21][30]~q ),
	.datac(\reg_file[29][30]~q ),
	.datad(\Mux1~0_combout ),
	.cin(gnd),
	.combout(\Mux1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~1 .lut_mask = 16'hF588;
defparam \Mux1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y29_N22
cycloneive_lcell_comb \Mux1~7 (
// Equation(s):
// \Mux1~7_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[27][30]~q )) # (!\prif.imemload_id [24] & ((\reg_file[19][30]~q )))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[27][30]~q ),
	.datac(\reg_file[19][30]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux1~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~7 .lut_mask = 16'hEE50;
defparam \Mux1~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y27_N10
cycloneive_lcell_comb \Mux1~8 (
// Equation(s):
// \Mux1~8_combout  = (\Mux1~7_combout  & (((\reg_file[31][30]~q ) # (!\prif.imemload_id [23])))) # (!\Mux1~7_combout  & (\reg_file[23][30]~q  & ((\prif.imemload_id [23]))))

	.dataa(\reg_file[23][30]~q ),
	.datab(\Mux1~7_combout ),
	.datac(\reg_file[31][30]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux1~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~8 .lut_mask = 16'hE2CC;
defparam \Mux1~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N6
cycloneive_lcell_comb \Mux1~3 (
// Equation(s):
// \Mux1~3_combout  = (\Mux1~2_combout  & (((\reg_file[30][30]~q )) # (!\prif.imemload_id [24]))) # (!\Mux1~2_combout  & (\prif.imemload_id [24] & (\reg_file[26][30]~q )))

	.dataa(\Mux1~2_combout ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[26][30]~q ),
	.datad(\reg_file[30][30]~q ),
	.cin(gnd),
	.combout(\Mux1~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~3 .lut_mask = 16'hEA62;
defparam \Mux1~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y33_N13
dffeas \reg_file[24][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~26_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[24][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[24][30] .is_wysiwyg = "true";
defparam \reg_file[24][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y33_N9
dffeas \reg_file[16][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][30] .is_wysiwyg = "true";
defparam \reg_file[16][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y33_N8
cycloneive_lcell_comb \Mux1~4 (
// Equation(s):
// \Mux1~4_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[20][30]~q ))) # (!\prif.imemload_id [23] & (\reg_file[16][30]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[16][30]~q ),
	.datad(\reg_file[20][30]~q ),
	.cin(gnd),
	.combout(\Mux1~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~4 .lut_mask = 16'hDC98;
defparam \Mux1~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y33_N12
cycloneive_lcell_comb \Mux1~5 (
// Equation(s):
// \Mux1~5_combout  = (\prif.imemload_id [24] & ((\Mux1~4_combout  & (\reg_file[28][30]~q )) # (!\Mux1~4_combout  & ((\reg_file[24][30]~q ))))) # (!\prif.imemload_id [24] & (((\Mux1~4_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[28][30]~q ),
	.datac(\reg_file[24][30]~q ),
	.datad(\Mux1~4_combout ),
	.cin(gnd),
	.combout(\Mux1~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~5 .lut_mask = 16'hDDA0;
defparam \Mux1~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N6
cycloneive_lcell_comb \Mux1~6 (
// Equation(s):
// \Mux1~6_combout  = (\prif.imemload_id [22] & ((\Mux1~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((!\prif.imemload_id [21] & \Mux1~5_combout ))))

	.dataa(\Mux1~3_combout ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux1~5_combout ),
	.cin(gnd),
	.combout(\Mux1~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~6 .lut_mask = 16'hCBC8;
defparam \Mux1~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y25_N12
cycloneive_lcell_comb \Mux1~17 (
// Equation(s):
// \Mux1~17_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[13][30]~q )) # (!\prif.imemload_id [21] & ((\reg_file[12][30]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[13][30]~q ),
	.datad(\reg_file[12][30]~q ),
	.cin(gnd),
	.combout(\Mux1~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~17 .lut_mask = 16'hD9C8;
defparam \Mux1~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N14
cycloneive_lcell_comb \Mux1~18 (
// Equation(s):
// \Mux1~18_combout  = (\prif.imemload_id [22] & ((\Mux1~17_combout  & (\reg_file[15][30]~q )) # (!\Mux1~17_combout  & ((\reg_file[14][30]~q ))))) # (!\prif.imemload_id [22] & (((\Mux1~17_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[15][30]~q ),
	.datac(\reg_file[14][30]~q ),
	.datad(\Mux1~17_combout ),
	.cin(gnd),
	.combout(\Mux1~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~18 .lut_mask = 16'hDDA0;
defparam \Mux1~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y30_N12
cycloneive_lcell_comb \reg_file[7][30]~feeder (
// Equation(s):
// \reg_file[7][30]~feeder_combout  = \reg_file_nxt[31][30]~70_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][30]~70_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[7][30]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[7][30]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[7][30]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X72_Y30_N13
dffeas \reg_file[7][30] (
	.clk(!CLK),
	.d(\reg_file[7][30]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~45_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[7][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[7][30] .is_wysiwyg = "true";
defparam \reg_file[7][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N8
cycloneive_lcell_comb \Mux1~10 (
// Equation(s):
// \Mux1~10_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[5][30]~q )) # (!\prif.imemload_id [21] & ((\reg_file[4][30]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[5][30]~q ),
	.datad(\reg_file[4][30]~q ),
	.cin(gnd),
	.combout(\Mux1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~10 .lut_mask = 16'hD9C8;
defparam \Mux1~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y27_N16
cycloneive_lcell_comb \Mux1~11 (
// Equation(s):
// \Mux1~11_combout  = (\prif.imemload_id [22] & ((\Mux1~10_combout  & (\reg_file[7][30]~q )) # (!\Mux1~10_combout  & ((\reg_file[6][30]~q ))))) # (!\prif.imemload_id [22] & (((\Mux1~10_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[7][30]~q ),
	.datac(\reg_file[6][30]~q ),
	.datad(\Mux1~10_combout ),
	.cin(gnd),
	.combout(\Mux1~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~11 .lut_mask = 16'hDDA0;
defparam \Mux1~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N18
cycloneive_lcell_comb \Mux1~13 (
// Equation(s):
// \Mux1~13_combout  = (\Mux1~12_combout  & (((\reg_file[11][30]~q )) # (!\prif.imemload_id [21]))) # (!\Mux1~12_combout  & (\prif.imemload_id [21] & ((\reg_file[9][30]~q ))))

	.dataa(\Mux1~12_combout ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[11][30]~q ),
	.datad(\reg_file[9][30]~q ),
	.cin(gnd),
	.combout(\Mux1~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~13 .lut_mask = 16'hE6A2;
defparam \Mux1~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y29_N3
dffeas \reg_file[1][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][30] .is_wysiwyg = "true";
defparam \reg_file[1][30] .power_up = "low";
// synopsys translate_on

// Location: FF_X67_Y29_N17
dffeas \reg_file[3][30] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][30]~70_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][30]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][30] .is_wysiwyg = "true";
defparam \reg_file[3][30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X67_Y29_N2
cycloneive_lcell_comb \Mux1~14 (
// Equation(s):
// \Mux1~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][30]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][30]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[1][30]~q ),
	.datad(\reg_file[3][30]~q ),
	.cin(gnd),
	.combout(\Mux1~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~14 .lut_mask = 16'hA820;
defparam \Mux1~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N2
cycloneive_lcell_comb \Mux1~15 (
// Equation(s):
// \Mux1~15_combout  = (\Mux1~14_combout ) # ((\reg_file[2][30]~q  & (\prif.imemload_id [22] & !\prif.imemload_id [21])))

	.dataa(\reg_file[2][30]~q ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux1~14_combout ),
	.cin(gnd),
	.combout(\Mux1~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~15 .lut_mask = 16'hFF08;
defparam \Mux1~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N16
cycloneive_lcell_comb \Mux1~16 (
// Equation(s):
// \Mux1~16_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\Mux1~13_combout )) # (!\prif.imemload_id [24] & ((\Mux1~15_combout )))))

	.dataa(\Mux1~13_combout ),
	.datab(prifimemload_id_23),
	.datac(prifimemload_id_24),
	.datad(\Mux1~15_combout ),
	.cin(gnd),
	.combout(\Mux1~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux1~16 .lut_mask = 16'hE3E0;
defparam \Mux1~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N16
cycloneive_lcell_comb \Mux2~3 (
// Equation(s):
// \Mux2~3_combout  = (\Mux2~2_combout  & ((\reg_file[30][29]~q ) # ((!\prif.imemload_id [23])))) # (!\Mux2~2_combout  & (((\reg_file[22][29]~q  & \prif.imemload_id [23]))))

	.dataa(\Mux2~2_combout ),
	.datab(\reg_file[30][29]~q ),
	.datac(\reg_file[22][29]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux2~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~3 .lut_mask = 16'hD8AA;
defparam \Mux2~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y31_N24
cycloneive_lcell_comb \reg_file[20][29]~feeder (
// Equation(s):
// \reg_file[20][29]~feeder_combout  = \reg_file_nxt[31][29]~71_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][29]~71_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[20][29]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[20][29]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[20][29]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X67_Y31_N25
dffeas \reg_file[20][29] (
	.clk(!CLK),
	.d(\reg_file[20][29]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][29] .is_wysiwyg = "true";
defparam \reg_file[20][29] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y32_N15
dffeas \reg_file[16][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][29] .is_wysiwyg = "true";
defparam \reg_file[16][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y32_N14
cycloneive_lcell_comb \Mux2~4 (
// Equation(s):
// \Mux2~4_combout  = (\prif.imemload_id [24] & ((\reg_file[24][29]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[16][29]~q  & !\prif.imemload_id [23]))))

	.dataa(\reg_file[24][29]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][29]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux2~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~4 .lut_mask = 16'hCCB8;
defparam \Mux2~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N14
cycloneive_lcell_comb \Mux2~5 (
// Equation(s):
// \Mux2~5_combout  = (\prif.imemload_id [23] & ((\Mux2~4_combout  & ((\reg_file[28][29]~q ))) # (!\Mux2~4_combout  & (\reg_file[20][29]~q )))) # (!\prif.imemload_id [23] & (((\Mux2~4_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[20][29]~q ),
	.datac(\reg_file[28][29]~q ),
	.datad(\Mux2~4_combout ),
	.cin(gnd),
	.combout(\Mux2~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~5 .lut_mask = 16'hF588;
defparam \Mux2~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N10
cycloneive_lcell_comb \Mux2~6 (
// Equation(s):
// \Mux2~6_combout  = (\prif.imemload_id [22] & ((\Mux2~3_combout ) # ((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (((!\prif.imemload_id [21] & \Mux2~5_combout ))))

	.dataa(\Mux2~3_combout ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux2~5_combout ),
	.cin(gnd),
	.combout(\Mux2~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~6 .lut_mask = 16'hCBC8;
defparam \Mux2~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N30
cycloneive_lcell_comb \Mux2~0 (
// Equation(s):
// \Mux2~0_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[21][29]~q ))) # (!\prif.imemload_id [23] & (\reg_file[17][29]~q ))))

	.dataa(\reg_file[17][29]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[21][29]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux2~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~0 .lut_mask = 16'hFC22;
defparam \Mux2~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y28_N2
cycloneive_lcell_comb \Mux2~1 (
// Equation(s):
// \Mux2~1_combout  = (\prif.imemload_id [24] & ((\Mux2~0_combout  & (\reg_file[29][29]~q )) # (!\Mux2~0_combout  & ((\reg_file[25][29]~q ))))) # (!\prif.imemload_id [24] & (((\Mux2~0_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[29][29]~q ),
	.datac(\Mux2~0_combout ),
	.datad(\reg_file[25][29]~q ),
	.cin(gnd),
	.combout(\Mux2~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~1 .lut_mask = 16'hDAD0;
defparam \Mux2~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N24
cycloneive_lcell_comb \Mux2~7 (
// Equation(s):
// \Mux2~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][29]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][29]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][29]~q ),
	.datad(\reg_file[23][29]~q ),
	.cin(gnd),
	.combout(\Mux2~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~7 .lut_mask = 16'hDC98;
defparam \Mux2~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y26_N18
cycloneive_lcell_comb \Mux2~8 (
// Equation(s):
// \Mux2~8_combout  = (\Mux2~7_combout  & (((\reg_file[31][29]~q ) # (!\prif.imemload_id [24])))) # (!\Mux2~7_combout  & (\reg_file[27][29]~q  & ((\prif.imemload_id [24]))))

	.dataa(\Mux2~7_combout ),
	.datab(\reg_file[27][29]~q ),
	.datac(\reg_file[31][29]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux2~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~8 .lut_mask = 16'hE4AA;
defparam \Mux2~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N16
cycloneive_lcell_comb \Mux2~12 (
// Equation(s):
// \Mux2~12_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[5][29]~q )) # (!\prif.imemload_id [21] & ((\reg_file[4][29]~q )))))

	.dataa(\reg_file[5][29]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[4][29]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux2~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~12 .lut_mask = 16'hEE30;
defparam \Mux2~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y28_N10
cycloneive_lcell_comb \Mux2~13 (
// Equation(s):
// \Mux2~13_combout  = (\prif.imemload_id [22] & ((\Mux2~12_combout  & (\reg_file[7][29]~q )) # (!\Mux2~12_combout  & ((\reg_file[6][29]~q ))))) # (!\prif.imemload_id [22] & (\Mux2~12_combout ))

	.dataa(prifimemload_id_22),
	.datab(\Mux2~12_combout ),
	.datac(\reg_file[7][29]~q ),
	.datad(\reg_file[6][29]~q ),
	.cin(gnd),
	.combout(\Mux2~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~13 .lut_mask = 16'hE6C4;
defparam \Mux2~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N14
cycloneive_lcell_comb \Mux2~14 (
// Equation(s):
// \Mux2~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][29]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][29]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[3][29]~q ),
	.datad(\reg_file[1][29]~q ),
	.cin(gnd),
	.combout(\Mux2~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~14 .lut_mask = 16'hC480;
defparam \Mux2~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y27_N22
cycloneive_lcell_comb \Mux2~15 (
// Equation(s):
// \Mux2~15_combout  = (\Mux2~14_combout ) # ((\reg_file[2][29]~q  & (\prif.imemload_id [22] & !\prif.imemload_id [21])))

	.dataa(\reg_file[2][29]~q ),
	.datab(prifimemload_id_22),
	.datac(\Mux2~14_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux2~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~15 .lut_mask = 16'hF0F8;
defparam \Mux2~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N30
cycloneive_lcell_comb \Mux2~16 (
// Equation(s):
// \Mux2~16_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\Mux2~13_combout )) # (!\prif.imemload_id [23] & ((\Mux2~15_combout )))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\Mux2~13_combout ),
	.datad(\Mux2~15_combout ),
	.cin(gnd),
	.combout(\Mux2~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~16 .lut_mask = 16'hD9C8;
defparam \Mux2~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N20
cycloneive_lcell_comb \Mux2~17 (
// Equation(s):
// \Mux2~17_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[13][29]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & ((\reg_file[12][29]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[13][29]~q ),
	.datad(\reg_file[12][29]~q ),
	.cin(gnd),
	.combout(\Mux2~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~17 .lut_mask = 16'hB9A8;
defparam \Mux2~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N4
cycloneive_lcell_comb \Mux2~18 (
// Equation(s):
// \Mux2~18_combout  = (\prif.imemload_id [22] & ((\Mux2~17_combout  & (\reg_file[15][29]~q )) # (!\Mux2~17_combout  & ((\reg_file[14][29]~q ))))) # (!\prif.imemload_id [22] & (\Mux2~17_combout ))

	.dataa(prifimemload_id_22),
	.datab(\Mux2~17_combout ),
	.datac(\reg_file[15][29]~q ),
	.datad(\reg_file[14][29]~q ),
	.cin(gnd),
	.combout(\Mux2~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~18 .lut_mask = 16'hE6C4;
defparam \Mux2~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X70_Y33_N9
dffeas \reg_file[9][29] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][29]~71_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~34_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[9][29]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[9][29] .is_wysiwyg = "true";
defparam \reg_file[9][29] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N18
cycloneive_lcell_comb \Mux2~10 (
// Equation(s):
// \Mux2~10_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[10][29]~q ))) # (!\prif.imemload_id [22] & (\reg_file[8][29]~q ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[8][29]~q ),
	.datad(\reg_file[10][29]~q ),
	.cin(gnd),
	.combout(\Mux2~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~10 .lut_mask = 16'hDC98;
defparam \Mux2~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y33_N8
cycloneive_lcell_comb \Mux2~11 (
// Equation(s):
// \Mux2~11_combout  = (\prif.imemload_id [21] & ((\Mux2~10_combout  & (\reg_file[11][29]~q )) # (!\Mux2~10_combout  & ((\reg_file[9][29]~q ))))) # (!\prif.imemload_id [21] & (((\Mux2~10_combout ))))

	.dataa(\reg_file[11][29]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[9][29]~q ),
	.datad(\Mux2~10_combout ),
	.cin(gnd),
	.combout(\Mux2~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux2~11 .lut_mask = 16'hBBC0;
defparam \Mux2~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N26
cycloneive_lcell_comb \Mux5~7 (
// Equation(s):
// \Mux5~7_combout  = (\prif.imemload_id [24] & ((\reg_file[27][26]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[19][26]~q  & !\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[27][26]~q ),
	.datac(\reg_file[19][26]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux5~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~7 .lut_mask = 16'hAAD8;
defparam \Mux5~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N12
cycloneive_lcell_comb \Mux5~8 (
// Equation(s):
// \Mux5~8_combout  = (\Mux5~7_combout  & (((\reg_file[31][26]~q )) # (!\prif.imemload_id [23]))) # (!\Mux5~7_combout  & (\prif.imemload_id [23] & ((\reg_file[23][26]~q ))))

	.dataa(\Mux5~7_combout ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[31][26]~q ),
	.datad(\reg_file[23][26]~q ),
	.cin(gnd),
	.combout(\Mux5~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~8 .lut_mask = 16'hE6A2;
defparam \Mux5~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N2
cycloneive_lcell_comb \Mux5~0 (
// Equation(s):
// \Mux5~0_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][26]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][26]~q )))))

	.dataa(\reg_file[25][26]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[17][26]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux5~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~0 .lut_mask = 16'hEE30;
defparam \Mux5~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y31_N10
cycloneive_lcell_comb \Mux5~1 (
// Equation(s):
// \Mux5~1_combout  = (\prif.imemload_id [23] & ((\Mux5~0_combout  & ((\reg_file[29][26]~q ))) # (!\Mux5~0_combout  & (\reg_file[21][26]~q )))) # (!\prif.imemload_id [23] & (((\Mux5~0_combout ))))

	.dataa(\reg_file[21][26]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[29][26]~q ),
	.datad(\Mux5~0_combout ),
	.cin(gnd),
	.combout(\Mux5~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~1 .lut_mask = 16'hF388;
defparam \Mux5~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y32_N11
dffeas \reg_file[16][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][26] .is_wysiwyg = "true";
defparam \reg_file[16][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N0
cycloneive_lcell_comb \Mux5~4 (
// Equation(s):
// \Mux5~4_combout  = (\prif.imemload_id [23] & (((\reg_file[20][26]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[16][26]~q  & ((!\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[16][26]~q ),
	.datac(\reg_file[20][26]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux5~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~4 .lut_mask = 16'hAAE4;
defparam \Mux5~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y32_N14
cycloneive_lcell_comb \Mux5~5 (
// Equation(s):
// \Mux5~5_combout  = (\Mux5~4_combout  & (((\reg_file[28][26]~q ) # (!\prif.imemload_id [24])))) # (!\Mux5~4_combout  & (\reg_file[24][26]~q  & ((\prif.imemload_id [24]))))

	.dataa(\reg_file[24][26]~q ),
	.datab(\Mux5~4_combout ),
	.datac(\reg_file[28][26]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux5~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~5 .lut_mask = 16'hE2CC;
defparam \Mux5~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y31_N29
dffeas \reg_file[18][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][26] .is_wysiwyg = "true";
defparam \reg_file[18][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y31_N28
cycloneive_lcell_comb \Mux5~2 (
// Equation(s):
// \Mux5~2_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & (\reg_file[22][26]~q )) # (!\prif.imemload_id [23] & ((\reg_file[18][26]~q )))))

	.dataa(\reg_file[22][26]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[18][26]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux5~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~2 .lut_mask = 16'hEE30;
defparam \Mux5~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X68_Y30_N21
dffeas \reg_file[26][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][26] .is_wysiwyg = "true";
defparam \reg_file[26][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N20
cycloneive_lcell_comb \Mux5~3 (
// Equation(s):
// \Mux5~3_combout  = (\prif.imemload_id [24] & ((\Mux5~2_combout  & (\reg_file[30][26]~q )) # (!\Mux5~2_combout  & ((\reg_file[26][26]~q ))))) # (!\prif.imemload_id [24] & (((\Mux5~2_combout ))))

	.dataa(\reg_file[30][26]~q ),
	.datab(prifimemload_id_24),
	.datac(\Mux5~2_combout ),
	.datad(\reg_file[26][26]~q ),
	.cin(gnd),
	.combout(\Mux5~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~3 .lut_mask = 16'hBCB0;
defparam \Mux5~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y34_N18
cycloneive_lcell_comb \Mux5~6 (
// Equation(s):
// \Mux5~6_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21]) # (\Mux5~3_combout )))) # (!\prif.imemload_id [22] & (\Mux5~5_combout  & (!\prif.imemload_id [21])))

	.dataa(\Mux5~5_combout ),
	.datab(prifimemload_id_22),
	.datac(prifimemload_id_21),
	.datad(\Mux5~3_combout ),
	.cin(gnd),
	.combout(\Mux5~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~6 .lut_mask = 16'hCEC2;
defparam \Mux5~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N11
dffeas \reg_file[12][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][26] .is_wysiwyg = "true";
defparam \reg_file[12][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N10
cycloneive_lcell_comb \Mux5~17 (
// Equation(s):
// \Mux5~17_combout  = (\prif.imemload_id [21] & ((\reg_file[13][26]~q ) # ((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (((\reg_file[12][26]~q  & !\prif.imemload_id [22]))))

	.dataa(\reg_file[13][26]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[12][26]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux5~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~17 .lut_mask = 16'hCCB8;
defparam \Mux5~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N2
cycloneive_lcell_comb \Mux5~18 (
// Equation(s):
// \Mux5~18_combout  = (\prif.imemload_id [22] & ((\Mux5~17_combout  & ((\reg_file[15][26]~q ))) # (!\Mux5~17_combout  & (\reg_file[14][26]~q )))) # (!\prif.imemload_id [22] & (((\Mux5~17_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[14][26]~q ),
	.datac(\reg_file[15][26]~q ),
	.datad(\Mux5~17_combout ),
	.cin(gnd),
	.combout(\Mux5~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~18 .lut_mask = 16'hF588;
defparam \Mux5~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y28_N31
dffeas \reg_file[4][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][26] .is_wysiwyg = "true";
defparam \reg_file[4][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N30
cycloneive_lcell_comb \Mux5~10 (
// Equation(s):
// \Mux5~10_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[5][26]~q )) # (!\prif.imemload_id [21] & ((\reg_file[4][26]~q )))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[5][26]~q ),
	.datac(\reg_file[4][26]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux5~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~10 .lut_mask = 16'hEE50;
defparam \Mux5~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N8
cycloneive_lcell_comb \Mux5~11 (
// Equation(s):
// \Mux5~11_combout  = (\Mux5~10_combout  & (((\reg_file[7][26]~q )) # (!\prif.imemload_id [22]))) # (!\Mux5~10_combout  & (\prif.imemload_id [22] & (\reg_file[6][26]~q )))

	.dataa(\Mux5~10_combout ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[6][26]~q ),
	.datad(\reg_file[7][26]~q ),
	.cin(gnd),
	.combout(\Mux5~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~11 .lut_mask = 16'hEA62;
defparam \Mux5~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y32_N6
cycloneive_lcell_comb \Mux5~14 (
// Equation(s):
// \Mux5~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][26]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][26]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][26]~q ),
	.datad(\reg_file[1][26]~q ),
	.cin(gnd),
	.combout(\Mux5~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~14 .lut_mask = 16'hA280;
defparam \Mux5~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N14
cycloneive_lcell_comb \Mux5~15 (
// Equation(s):
// \Mux5~15_combout  = (\Mux5~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][26]~q  & !\prif.imemload_id [21])))

	.dataa(prifimemload_id_22),
	.datab(\Mux5~14_combout ),
	.datac(\reg_file[2][26]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux5~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~15 .lut_mask = 16'hCCEC;
defparam \Mux5~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N23
dffeas \reg_file[8][26] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][26]~91_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][26]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][26] .is_wysiwyg = "true";
defparam \reg_file[8][26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N22
cycloneive_lcell_comb \Mux5~12 (
// Equation(s):
// \Mux5~12_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[10][26]~q )) # (!\prif.imemload_id [22] & ((\reg_file[8][26]~q )))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[10][26]~q ),
	.datac(\reg_file[8][26]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux5~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~12 .lut_mask = 16'hEE50;
defparam \Mux5~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N22
cycloneive_lcell_comb \Mux5~13 (
// Equation(s):
// \Mux5~13_combout  = (\prif.imemload_id [21] & ((\Mux5~12_combout  & (\reg_file[11][26]~q )) # (!\Mux5~12_combout  & ((\reg_file[9][26]~q ))))) # (!\prif.imemload_id [21] & (((\Mux5~12_combout ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[11][26]~q ),
	.datac(\reg_file[9][26]~q ),
	.datad(\Mux5~12_combout ),
	.cin(gnd),
	.combout(\Mux5~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~13 .lut_mask = 16'hDDA0;
defparam \Mux5~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N20
cycloneive_lcell_comb \Mux5~16 (
// Equation(s):
// \Mux5~16_combout  = (\prif.imemload_id [24] & (((\Mux5~13_combout ) # (\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (\Mux5~15_combout  & ((!\prif.imemload_id [23]))))

	.dataa(prifimemload_id_24),
	.datab(\Mux5~15_combout ),
	.datac(\Mux5~13_combout ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux5~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux5~16 .lut_mask = 16'hAAE4;
defparam \Mux5~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N16
cycloneive_lcell_comb \Mux6~0 (
// Equation(s):
// \Mux6~0_combout  = (\prif.imemload_id [24] & (((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[21][25]~q ))) # (!\prif.imemload_id [23] & (\reg_file[17][25]~q ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[17][25]~q ),
	.datac(prifimemload_id_23),
	.datad(\reg_file[21][25]~q ),
	.cin(gnd),
	.combout(\Mux6~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~0 .lut_mask = 16'hF4A4;
defparam \Mux6~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y29_N2
cycloneive_lcell_comb \Mux6~1 (
// Equation(s):
// \Mux6~1_combout  = (\prif.imemload_id [24] & ((\Mux6~0_combout  & ((\reg_file[29][25]~q ))) # (!\Mux6~0_combout  & (\reg_file[25][25]~q )))) # (!\prif.imemload_id [24] & (((\Mux6~0_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[25][25]~q ),
	.datac(\reg_file[29][25]~q ),
	.datad(\Mux6~0_combout ),
	.cin(gnd),
	.combout(\Mux6~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~1 .lut_mask = 16'hF588;
defparam \Mux6~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N20
cycloneive_lcell_comb \Mux6~7 (
// Equation(s):
// \Mux6~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][25]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][25]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][25]~q ),
	.datad(\reg_file[23][25]~q ),
	.cin(gnd),
	.combout(\Mux6~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~7 .lut_mask = 16'hDC98;
defparam \Mux6~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N12
cycloneive_lcell_comb \Mux6~8 (
// Equation(s):
// \Mux6~8_combout  = (\prif.imemload_id [24] & ((\Mux6~7_combout  & (\reg_file[31][25]~q )) # (!\Mux6~7_combout  & ((\reg_file[27][25]~q ))))) # (!\prif.imemload_id [24] & (((\Mux6~7_combout ))))

	.dataa(prifimemload_id_24),
	.datab(\reg_file[31][25]~q ),
	.datac(\reg_file[27][25]~q ),
	.datad(\Mux6~7_combout ),
	.cin(gnd),
	.combout(\Mux6~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~8 .lut_mask = 16'hDDA0;
defparam \Mux6~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N13
dffeas \reg_file[20][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~27_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[20][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[20][25] .is_wysiwyg = "true";
defparam \reg_file[20][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X66_Y35_N3
dffeas \reg_file[16][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][25] .is_wysiwyg = "true";
defparam \reg_file[16][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N2
cycloneive_lcell_comb \Mux6~4 (
// Equation(s):
// \Mux6~4_combout  = (\prif.imemload_id [24] & ((\reg_file[24][25]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[16][25]~q  & !\prif.imemload_id [23]))))

	.dataa(\reg_file[24][25]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][25]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux6~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~4 .lut_mask = 16'hCCB8;
defparam \Mux6~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y34_N24
cycloneive_lcell_comb \Mux6~5 (
// Equation(s):
// \Mux6~5_combout  = (\prif.imemload_id [23] & ((\Mux6~4_combout  & ((\reg_file[28][25]~q ))) # (!\Mux6~4_combout  & (\reg_file[20][25]~q )))) # (!\prif.imemload_id [23] & (((\Mux6~4_combout ))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[20][25]~q ),
	.datac(\reg_file[28][25]~q ),
	.datad(\Mux6~4_combout ),
	.cin(gnd),
	.combout(\Mux6~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~5 .lut_mask = 16'hF588;
defparam \Mux6~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N8
cycloneive_lcell_comb \Mux6~3 (
// Equation(s):
// \Mux6~3_combout  = (\Mux6~2_combout  & ((\reg_file[30][25]~q ) # ((!\prif.imemload_id [23])))) # (!\Mux6~2_combout  & (((\prif.imemload_id [23] & \reg_file[22][25]~q ))))

	.dataa(\Mux6~2_combout ),
	.datab(\reg_file[30][25]~q ),
	.datac(prifimemload_id_23),
	.datad(\reg_file[22][25]~q ),
	.cin(gnd),
	.combout(\Mux6~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~3 .lut_mask = 16'hDA8A;
defparam \Mux6~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y30_N10
cycloneive_lcell_comb \Mux6~6 (
// Equation(s):
// \Mux6~6_combout  = (\prif.imemload_id [22] & (((\Mux6~3_combout ) # (\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (\Mux6~5_combout  & ((!\prif.imemload_id [21]))))

	.dataa(\Mux6~5_combout ),
	.datab(prifimemload_id_22),
	.datac(\Mux6~3_combout ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux6~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~6 .lut_mask = 16'hCCE2;
defparam \Mux6~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y25_N28
cycloneive_lcell_comb \Mux6~10 (
// Equation(s):
// \Mux6~10_combout  = (\prif.imemload_id [22] & (((\reg_file[10][25]~q ) # (\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & (\reg_file[8][25]~q  & ((!\prif.imemload_id [21]))))

	.dataa(\reg_file[8][25]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[10][25]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux6~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~10 .lut_mask = 16'hCCE2;
defparam \Mux6~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y25_N24
cycloneive_lcell_comb \Mux6~11 (
// Equation(s):
// \Mux6~11_combout  = (\prif.imemload_id [21] & ((\Mux6~10_combout  & (\reg_file[11][25]~q )) # (!\Mux6~10_combout  & ((\reg_file[9][25]~q ))))) # (!\prif.imemload_id [21] & (((\Mux6~10_combout ))))

	.dataa(\reg_file[11][25]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[9][25]~q ),
	.datad(\Mux6~10_combout ),
	.cin(gnd),
	.combout(\Mux6~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~11 .lut_mask = 16'hBBC0;
defparam \Mux6~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y29_N17
dffeas \reg_file[3][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~46_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[3][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[3][25] .is_wysiwyg = "true";
defparam \reg_file[3][25] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y29_N3
dffeas \reg_file[1][25] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][25]~95_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~47_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[1][25]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[1][25] .is_wysiwyg = "true";
defparam \reg_file[1][25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y29_N16
cycloneive_lcell_comb \Mux6~14 (
// Equation(s):
// \Mux6~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[3][25]~q )) # (!\prif.imemload_id [22] & ((\reg_file[1][25]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[3][25]~q ),
	.datad(\reg_file[1][25]~q ),
	.cin(gnd),
	.combout(\Mux6~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~14 .lut_mask = 16'hA280;
defparam \Mux6~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N8
cycloneive_lcell_comb \Mux6~15 (
// Equation(s):
// \Mux6~15_combout  = (\Mux6~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][25]~q  & !\prif.imemload_id [21])))

	.dataa(prifimemload_id_22),
	.datab(\Mux6~14_combout ),
	.datac(\reg_file[2][25]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux6~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~15 .lut_mask = 16'hCCEC;
defparam \Mux6~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N6
cycloneive_lcell_comb \Mux6~12 (
// Equation(s):
// \Mux6~12_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[5][25]~q ))) # (!\prif.imemload_id [21] & (\reg_file[4][25]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[4][25]~q ),
	.datad(\reg_file[5][25]~q ),
	.cin(gnd),
	.combout(\Mux6~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~12 .lut_mask = 16'hDC98;
defparam \Mux6~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N2
cycloneive_lcell_comb \Mux6~13 (
// Equation(s):
// \Mux6~13_combout  = (\prif.imemload_id [22] & ((\Mux6~12_combout  & ((\reg_file[7][25]~q ))) # (!\Mux6~12_combout  & (\reg_file[6][25]~q )))) # (!\prif.imemload_id [22] & (((\Mux6~12_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[6][25]~q ),
	.datac(\reg_file[7][25]~q ),
	.datad(\Mux6~12_combout ),
	.cin(gnd),
	.combout(\Mux6~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~13 .lut_mask = 16'hF588;
defparam \Mux6~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N26
cycloneive_lcell_comb \Mux6~16 (
// Equation(s):
// \Mux6~16_combout  = (\prif.imemload_id [23] & ((\prif.imemload_id [24]) # ((\Mux6~13_combout )))) # (!\prif.imemload_id [23] & (!\prif.imemload_id [24] & (\Mux6~15_combout )))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\Mux6~15_combout ),
	.datad(\Mux6~13_combout ),
	.cin(gnd),
	.combout(\Mux6~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~16 .lut_mask = 16'hBA98;
defparam \Mux6~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X62_Y26_N18
cycloneive_lcell_comb \Mux6~17 (
// Equation(s):
// \Mux6~17_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22]) # ((\reg_file[13][25]~q )))) # (!\prif.imemload_id [21] & (!\prif.imemload_id [22] & (\reg_file[12][25]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[12][25]~q ),
	.datad(\reg_file[13][25]~q ),
	.cin(gnd),
	.combout(\Mux6~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~17 .lut_mask = 16'hBA98;
defparam \Mux6~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y26_N26
cycloneive_lcell_comb \Mux6~18 (
// Equation(s):
// \Mux6~18_combout  = (\prif.imemload_id [22] & ((\Mux6~17_combout  & ((\reg_file[15][25]~q ))) # (!\Mux6~17_combout  & (\reg_file[14][25]~q )))) # (!\prif.imemload_id [22] & (((\Mux6~17_combout ))))

	.dataa(\reg_file[14][25]~q ),
	.datab(\reg_file[15][25]~q ),
	.datac(prifimemload_id_22),
	.datad(\Mux6~17_combout ),
	.cin(gnd),
	.combout(\Mux6~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux6~18 .lut_mask = 16'hCFA0;
defparam \Mux6~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N14
cycloneive_lcell_comb \Mux3~7 (
// Equation(s):
// \Mux3~7_combout  = (\prif.imemload_id [24] & ((\prif.imemload_id [23]) # ((\reg_file[27][28]~q )))) # (!\prif.imemload_id [24] & (!\prif.imemload_id [23] & (\reg_file[19][28]~q )))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][28]~q ),
	.datad(\reg_file[27][28]~q ),
	.cin(gnd),
	.combout(\Mux3~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~7 .lut_mask = 16'hBA98;
defparam \Mux3~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N0
cycloneive_lcell_comb \Mux3~8 (
// Equation(s):
// \Mux3~8_combout  = (\prif.imemload_id [23] & ((\Mux3~7_combout  & (\reg_file[31][28]~q )) # (!\Mux3~7_combout  & ((\reg_file[23][28]~q ))))) # (!\prif.imemload_id [23] & (\Mux3~7_combout ))

	.dataa(prifimemload_id_23),
	.datab(\Mux3~7_combout ),
	.datac(\reg_file[31][28]~q ),
	.datad(\reg_file[23][28]~q ),
	.cin(gnd),
	.combout(\Mux3~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~8 .lut_mask = 16'hE6C4;
defparam \Mux3~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N0
cycloneive_lcell_comb \Mux3~0 (
// Equation(s):
// \Mux3~0_combout  = (\prif.imemload_id [23] & (((\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[25][28]~q )) # (!\prif.imemload_id [24] & ((\reg_file[17][28]~q )))))

	.dataa(\reg_file[25][28]~q ),
	.datab(prifimemload_id_23),
	.datac(\reg_file[17][28]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux3~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~0 .lut_mask = 16'hEE30;
defparam \Mux3~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y30_N6
cycloneive_lcell_comb \Mux3~1 (
// Equation(s):
// \Mux3~1_combout  = (\Mux3~0_combout  & (((\reg_file[29][28]~q ) # (!\prif.imemload_id [23])))) # (!\Mux3~0_combout  & (\reg_file[21][28]~q  & ((\prif.imemload_id [23]))))

	.dataa(\reg_file[21][28]~q ),
	.datab(\Mux3~0_combout ),
	.datac(\reg_file[29][28]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux3~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~1 .lut_mask = 16'hE2CC;
defparam \Mux3~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y33_N18
cycloneive_lcell_comb \Mux3~5 (
// Equation(s):
// \Mux3~5_combout  = (\Mux3~4_combout  & (((\reg_file[28][28]~q ) # (!\prif.imemload_id [24])))) # (!\Mux3~4_combout  & (\reg_file[24][28]~q  & ((\prif.imemload_id [24]))))

	.dataa(\Mux3~4_combout ),
	.datab(\reg_file[24][28]~q ),
	.datac(\reg_file[28][28]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux3~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~5 .lut_mask = 16'hE4AA;
defparam \Mux3~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N9
dffeas \reg_file[26][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~21_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[26][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[26][28] .is_wysiwyg = "true";
defparam \reg_file[26][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y31_N14
cycloneive_lcell_comb \Mux3~3 (
// Equation(s):
// \Mux3~3_combout  = (\Mux3~2_combout  & (((\reg_file[30][28]~q )) # (!\prif.imemload_id [24]))) # (!\Mux3~2_combout  & (\prif.imemload_id [24] & ((\reg_file[26][28]~q ))))

	.dataa(\Mux3~2_combout ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[30][28]~q ),
	.datad(\reg_file[26][28]~q ),
	.cin(gnd),
	.combout(\Mux3~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~3 .lut_mask = 16'hE6A2;
defparam \Mux3~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y34_N14
cycloneive_lcell_comb \Mux3~6 (
// Equation(s):
// \Mux3~6_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\Mux3~3_combout ))) # (!\prif.imemload_id [22] & (\Mux3~5_combout ))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux3~5_combout ),
	.datad(\Mux3~3_combout ),
	.cin(gnd),
	.combout(\Mux3~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~6 .lut_mask = 16'hDC98;
defparam \Mux3~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y28_N27
dffeas \reg_file[5][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[5][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[5][28] .is_wysiwyg = "true";
defparam \reg_file[5][28] .power_up = "low";
// synopsys translate_on

// Location: FF_X73_Y28_N13
dffeas \reg_file[4][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~44_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[4][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[4][28] .is_wysiwyg = "true";
defparam \reg_file[4][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N26
cycloneive_lcell_comb \Mux3~10 (
// Equation(s):
// \Mux3~10_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[5][28]~q )) # (!\prif.imemload_id [21] & ((\reg_file[4][28]~q )))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[5][28]~q ),
	.datad(\reg_file[4][28]~q ),
	.cin(gnd),
	.combout(\Mux3~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~10 .lut_mask = 16'hD9C8;
defparam \Mux3~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y28_N18
cycloneive_lcell_comb \Mux3~11 (
// Equation(s):
// \Mux3~11_combout  = (\prif.imemload_id [22] & ((\Mux3~10_combout  & (\reg_file[7][28]~q )) # (!\Mux3~10_combout  & ((\reg_file[6][28]~q ))))) # (!\prif.imemload_id [22] & (((\Mux3~10_combout ))))

	.dataa(\reg_file[7][28]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[6][28]~q ),
	.datad(\Mux3~10_combout ),
	.cin(gnd),
	.combout(\Mux3~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~11 .lut_mask = 16'hBBC0;
defparam \Mux3~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N22
cycloneive_lcell_comb \Mux3~14 (
// Equation(s):
// \Mux3~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][28]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][28]~q ))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[1][28]~q ),
	.datac(prifimemload_id_22),
	.datad(\reg_file[3][28]~q ),
	.cin(gnd),
	.combout(\Mux3~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~14 .lut_mask = 16'hA808;
defparam \Mux3~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N10
cycloneive_lcell_comb \Mux3~15 (
// Equation(s):
// \Mux3~15_combout  = (\Mux3~14_combout ) # ((\prif.imemload_id [22] & (\reg_file[2][28]~q  & !\prif.imemload_id [21])))

	.dataa(prifimemload_id_22),
	.datab(\Mux3~14_combout ),
	.datac(\reg_file[2][28]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux3~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~15 .lut_mask = 16'hCCEC;
defparam \Mux3~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X69_Y35_N31
dffeas \reg_file[8][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~36_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[8][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[8][28] .is_wysiwyg = "true";
defparam \reg_file[8][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N30
cycloneive_lcell_comb \Mux3~12 (
// Equation(s):
// \Mux3~12_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[10][28]~q )) # (!\prif.imemload_id [22] & ((\reg_file[8][28]~q )))))

	.dataa(prifimemload_id_21),
	.datab(\reg_file[10][28]~q ),
	.datac(\reg_file[8][28]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux3~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~12 .lut_mask = 16'hEE50;
defparam \Mux3~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N0
cycloneive_lcell_comb \Mux3~13 (
// Equation(s):
// \Mux3~13_combout  = (\Mux3~12_combout  & ((\reg_file[11][28]~q ) # ((!\prif.imemload_id [21])))) # (!\Mux3~12_combout  & (((\reg_file[9][28]~q  & \prif.imemload_id [21]))))

	.dataa(\reg_file[11][28]~q ),
	.datab(\Mux3~12_combout ),
	.datac(\reg_file[9][28]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux3~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~13 .lut_mask = 16'hB8CC;
defparam \Mux3~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y34_N4
cycloneive_lcell_comb \Mux3~16 (
// Equation(s):
// \Mux3~16_combout  = (\prif.imemload_id [24] & (((\Mux3~13_combout ) # (\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (\Mux3~15_combout  & ((!\prif.imemload_id [23]))))

	.dataa(\Mux3~15_combout ),
	.datab(\Mux3~13_combout ),
	.datac(prifimemload_id_24),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux3~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~16 .lut_mask = 16'hF0CA;
defparam \Mux3~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X73_Y32_N31
dffeas \reg_file[12][28] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][28]~90_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~40_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[12][28]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[12][28] .is_wysiwyg = "true";
defparam \reg_file[12][28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N30
cycloneive_lcell_comb \Mux3~17 (
// Equation(s):
// \Mux3~17_combout  = (\prif.imemload_id [22] & (\prif.imemload_id [21])) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & ((\reg_file[13][28]~q ))) # (!\prif.imemload_id [21] & (\reg_file[12][28]~q ))))

	.dataa(prifimemload_id_22),
	.datab(prifimemload_id_21),
	.datac(\reg_file[12][28]~q ),
	.datad(\reg_file[13][28]~q ),
	.cin(gnd),
	.combout(\Mux3~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~17 .lut_mask = 16'hDC98;
defparam \Mux3~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y31_N22
cycloneive_lcell_comb \Mux3~18 (
// Equation(s):
// \Mux3~18_combout  = (\prif.imemload_id [22] & ((\Mux3~17_combout  & (\reg_file[15][28]~q )) # (!\Mux3~17_combout  & ((\reg_file[14][28]~q ))))) # (!\prif.imemload_id [22] & (((\Mux3~17_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[15][28]~q ),
	.datac(\Mux3~17_combout ),
	.datad(\reg_file[14][28]~q ),
	.cin(gnd),
	.combout(\Mux3~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux3~18 .lut_mask = 16'hDAD0;
defparam \Mux3~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X67_Y32_N12
cycloneive_lcell_comb \Mux4~0 (
// Equation(s):
// \Mux4~0_combout  = (\prif.imemload_id [23] & (((\reg_file[21][27]~q ) # (\prif.imemload_id [24])))) # (!\prif.imemload_id [23] & (\reg_file[17][27]~q  & ((!\prif.imemload_id [24]))))

	.dataa(prifimemload_id_23),
	.datab(\reg_file[17][27]~q ),
	.datac(\reg_file[21][27]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux4~0_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~0 .lut_mask = 16'hAAE4;
defparam \Mux4~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N0
cycloneive_lcell_comb \reg_file[25][27]~feeder (
// Equation(s):
// \reg_file[25][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][27]~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[25][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[25][27]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[25][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y28_N1
dffeas \reg_file[25][27] (
	.clk(!CLK),
	.d(\reg_file[25][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~17_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[25][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[25][27] .is_wysiwyg = "true";
defparam \reg_file[25][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N14
cycloneive_lcell_comb \Mux4~1 (
// Equation(s):
// \Mux4~1_combout  = (\Mux4~0_combout  & ((\reg_file[29][27]~q ) # ((!\prif.imemload_id [24])))) # (!\Mux4~0_combout  & (((\prif.imemload_id [24] & \reg_file[25][27]~q ))))

	.dataa(\reg_file[29][27]~q ),
	.datab(\Mux4~0_combout ),
	.datac(prifimemload_id_24),
	.datad(\reg_file[25][27]~q ),
	.cin(gnd),
	.combout(\Mux4~1_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~1 .lut_mask = 16'hBC8C;
defparam \Mux4~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y31_N12
cycloneive_lcell_comb \reg_file[18][27]~feeder (
// Equation(s):
// \reg_file[18][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(\reg_file_nxt[31][27]~81_combout ),
	.cin(gnd),
	.combout(\reg_file[18][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[18][27]~feeder .lut_mask = 16'hFF00;
defparam \reg_file[18][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X65_Y31_N13
dffeas \reg_file[18][27] (
	.clk(!CLK),
	.d(\reg_file[18][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~24_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[18][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[18][27] .is_wysiwyg = "true";
defparam \reg_file[18][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y28_N10
cycloneive_lcell_comb \Mux4~2 (
// Equation(s):
// \Mux4~2_combout  = (\prif.imemload_id [23] & (\prif.imemload_id [24])) # (!\prif.imemload_id [23] & ((\prif.imemload_id [24] & (\reg_file[26][27]~q )) # (!\prif.imemload_id [24] & ((\reg_file[18][27]~q )))))

	.dataa(prifimemload_id_23),
	.datab(prifimemload_id_24),
	.datac(\reg_file[26][27]~q ),
	.datad(\reg_file[18][27]~q ),
	.cin(gnd),
	.combout(\Mux4~2_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~2 .lut_mask = 16'hD9C8;
defparam \Mux4~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N4
cycloneive_lcell_comb \reg_file[22][27]~feeder (
// Equation(s):
// \reg_file[22][27]~feeder_combout  = \reg_file_nxt[31][27]~81_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(\reg_file_nxt[31][27]~81_combout ),
	.datad(gnd),
	.cin(gnd),
	.combout(\reg_file[22][27]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \reg_file[22][27]~feeder .lut_mask = 16'hF0F0;
defparam \reg_file[22][27]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X63_Y30_N5
dffeas \reg_file[22][27] (
	.clk(!CLK),
	.d(\reg_file[22][27]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\Decoder0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[22][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[22][27] .is_wysiwyg = "true";
defparam \reg_file[22][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X63_Y30_N22
cycloneive_lcell_comb \Mux4~3 (
// Equation(s):
// \Mux4~3_combout  = (\prif.imemload_id [23] & ((\Mux4~2_combout  & (\reg_file[30][27]~q )) # (!\Mux4~2_combout  & ((\reg_file[22][27]~q ))))) # (!\prif.imemload_id [23] & (\Mux4~2_combout ))

	.dataa(prifimemload_id_23),
	.datab(\Mux4~2_combout ),
	.datac(\reg_file[30][27]~q ),
	.datad(\reg_file[22][27]~q ),
	.cin(gnd),
	.combout(\Mux4~3_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~3 .lut_mask = 16'hE6C4;
defparam \Mux4~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X66_Y35_N31
dffeas \reg_file[16][27] (
	.clk(!CLK),
	.d(gnd),
	.asdata(\reg_file_nxt[31][27]~81_combout ),
	.clrn(nRST),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\Decoder0~28_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\reg_file[16][27]~q ),
	.prn(vcc));
// synopsys translate_off
defparam \reg_file[16][27] .is_wysiwyg = "true";
defparam \reg_file[16][27] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X66_Y35_N30
cycloneive_lcell_comb \Mux4~4 (
// Equation(s):
// \Mux4~4_combout  = (\prif.imemload_id [24] & ((\reg_file[24][27]~q ) # ((\prif.imemload_id [23])))) # (!\prif.imemload_id [24] & (((\reg_file[16][27]~q  & !\prif.imemload_id [23]))))

	.dataa(\reg_file[24][27]~q ),
	.datab(prifimemload_id_24),
	.datac(\reg_file[16][27]~q ),
	.datad(prifimemload_id_23),
	.cin(gnd),
	.combout(\Mux4~4_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~4 .lut_mask = 16'hCCB8;
defparam \Mux4~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y34_N6
cycloneive_lcell_comb \Mux4~5 (
// Equation(s):
// \Mux4~5_combout  = (\prif.imemload_id [23] & ((\Mux4~4_combout  & ((\reg_file[28][27]~q ))) # (!\Mux4~4_combout  & (\reg_file[20][27]~q )))) # (!\prif.imemload_id [23] & (((\Mux4~4_combout ))))

	.dataa(\reg_file[20][27]~q ),
	.datab(prifimemload_id_23),
	.datac(\Mux4~4_combout ),
	.datad(\reg_file[28][27]~q ),
	.cin(gnd),
	.combout(\Mux4~5_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~5 .lut_mask = 16'hF838;
defparam \Mux4~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N4
cycloneive_lcell_comb \Mux4~6 (
// Equation(s):
// \Mux4~6_combout  = (\prif.imemload_id [21] & (((\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\Mux4~3_combout )) # (!\prif.imemload_id [22] & ((\Mux4~5_combout )))))

	.dataa(prifimemload_id_21),
	.datab(\Mux4~3_combout ),
	.datac(prifimemload_id_22),
	.datad(\Mux4~5_combout ),
	.cin(gnd),
	.combout(\Mux4~6_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~6 .lut_mask = 16'hE5E0;
defparam \Mux4~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X70_Y27_N28
cycloneive_lcell_comb \Mux4~7 (
// Equation(s):
// \Mux4~7_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\reg_file[23][27]~q ))) # (!\prif.imemload_id [23] & (\reg_file[19][27]~q ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\reg_file[19][27]~q ),
	.datad(\reg_file[23][27]~q ),
	.cin(gnd),
	.combout(\Mux4~7_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~7 .lut_mask = 16'hDC98;
defparam \Mux4~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N6
cycloneive_lcell_comb \Mux4~8 (
// Equation(s):
// \Mux4~8_combout  = (\Mux4~7_combout  & (((\reg_file[31][27]~q ) # (!\prif.imemload_id [24])))) # (!\Mux4~7_combout  & (\reg_file[27][27]~q  & ((\prif.imemload_id [24]))))

	.dataa(\reg_file[27][27]~q ),
	.datab(\Mux4~7_combout ),
	.datac(\reg_file[31][27]~q ),
	.datad(prifimemload_id_24),
	.cin(gnd),
	.combout(\Mux4~8_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~8 .lut_mask = 16'hE2CC;
defparam \Mux4~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X69_Y35_N24
cycloneive_lcell_comb \Mux4~10 (
// Equation(s):
// \Mux4~10_combout  = (\prif.imemload_id [21] & (\prif.imemload_id [22])) # (!\prif.imemload_id [21] & ((\prif.imemload_id [22] & (\reg_file[10][27]~q )) # (!\prif.imemload_id [22] & ((\reg_file[8][27]~q )))))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\reg_file[10][27]~q ),
	.datad(\reg_file[8][27]~q ),
	.cin(gnd),
	.combout(\Mux4~10_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~10 .lut_mask = 16'hD9C8;
defparam \Mux4~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X68_Y35_N0
cycloneive_lcell_comb \Mux4~11 (
// Equation(s):
// \Mux4~11_combout  = (\Mux4~10_combout  & ((\reg_file[11][27]~q ) # ((!\prif.imemload_id [21])))) # (!\Mux4~10_combout  & (((\reg_file[9][27]~q  & \prif.imemload_id [21]))))

	.dataa(\reg_file[11][27]~q ),
	.datab(\Mux4~10_combout ),
	.datac(\reg_file[9][27]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux4~11_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~11 .lut_mask = 16'hB8CC;
defparam \Mux4~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N26
cycloneive_lcell_comb \Mux4~14 (
// Equation(s):
// \Mux4~14_combout  = (\prif.imemload_id [21] & ((\prif.imemload_id [22] & ((\reg_file[3][27]~q ))) # (!\prif.imemload_id [22] & (\reg_file[1][27]~q ))))

	.dataa(\reg_file[1][27]~q ),
	.datab(\reg_file[3][27]~q ),
	.datac(prifimemload_id_22),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux4~14_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~14 .lut_mask = 16'hCA00;
defparam \Mux4~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N0
cycloneive_lcell_comb \Mux4~15 (
// Equation(s):
// \Mux4~15_combout  = (\Mux4~14_combout ) # ((!\prif.imemload_id [21] & (\prif.imemload_id [22] & \reg_file[2][27]~q )))

	.dataa(prifimemload_id_21),
	.datab(prifimemload_id_22),
	.datac(\Mux4~14_combout ),
	.datad(\reg_file[2][27]~q ),
	.cin(gnd),
	.combout(\Mux4~15_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~15 .lut_mask = 16'hF4F0;
defparam \Mux4~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y28_N0
cycloneive_lcell_comb \Mux4~12 (
// Equation(s):
// \Mux4~12_combout  = (\prif.imemload_id [22] & (((\prif.imemload_id [21])))) # (!\prif.imemload_id [22] & ((\prif.imemload_id [21] & (\reg_file[5][27]~q )) # (!\prif.imemload_id [21] & ((\reg_file[4][27]~q )))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[5][27]~q ),
	.datac(\reg_file[4][27]~q ),
	.datad(prifimemload_id_21),
	.cin(gnd),
	.combout(\Mux4~12_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~12 .lut_mask = 16'hEE50;
defparam \Mux4~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X72_Y29_N2
cycloneive_lcell_comb \Mux4~13 (
// Equation(s):
// \Mux4~13_combout  = (\prif.imemload_id [22] & ((\Mux4~12_combout  & ((\reg_file[7][27]~q ))) # (!\Mux4~12_combout  & (\reg_file[6][27]~q )))) # (!\prif.imemload_id [22] & (((\Mux4~12_combout ))))

	.dataa(\reg_file[6][27]~q ),
	.datab(prifimemload_id_22),
	.datac(\reg_file[7][27]~q ),
	.datad(\Mux4~12_combout ),
	.cin(gnd),
	.combout(\Mux4~13_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~13 .lut_mask = 16'hF388;
defparam \Mux4~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X63_Y34_N18
cycloneive_lcell_comb \Mux4~16 (
// Equation(s):
// \Mux4~16_combout  = (\prif.imemload_id [24] & (\prif.imemload_id [23])) # (!\prif.imemload_id [24] & ((\prif.imemload_id [23] & ((\Mux4~13_combout ))) # (!\prif.imemload_id [23] & (\Mux4~15_combout ))))

	.dataa(prifimemload_id_24),
	.datab(prifimemload_id_23),
	.datac(\Mux4~15_combout ),
	.datad(\Mux4~13_combout ),
	.cin(gnd),
	.combout(\Mux4~16_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~16 .lut_mask = 16'hDC98;
defparam \Mux4~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X73_Y32_N4
cycloneive_lcell_comb \Mux4~17 (
// Equation(s):
// \Mux4~17_combout  = (\prif.imemload_id [21] & (((\reg_file[13][27]~q ) # (\prif.imemload_id [22])))) # (!\prif.imemload_id [21] & (\reg_file[12][27]~q  & ((!\prif.imemload_id [22]))))

	.dataa(\reg_file[12][27]~q ),
	.datab(prifimemload_id_21),
	.datac(\reg_file[13][27]~q ),
	.datad(prifimemload_id_22),
	.cin(gnd),
	.combout(\Mux4~17_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~17 .lut_mask = 16'hCCE2;
defparam \Mux4~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X65_Y29_N30
cycloneive_lcell_comb \Mux4~18 (
// Equation(s):
// \Mux4~18_combout  = (\prif.imemload_id [22] & ((\Mux4~17_combout  & ((\reg_file[15][27]~q ))) # (!\Mux4~17_combout  & (\reg_file[14][27]~q )))) # (!\prif.imemload_id [22] & (((\Mux4~17_combout ))))

	.dataa(prifimemload_id_22),
	.datab(\reg_file[14][27]~q ),
	.datac(\reg_file[15][27]~q ),
	.datad(\Mux4~17_combout ),
	.cin(gnd),
	.combout(\Mux4~18_combout ),
	.cout());
// synopsys translate_off
defparam \Mux4~18 .lut_mask = 16'hF588;
defparam \Mux4~18 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module memory_control (
	prifdmemren,
	prifdmemwen,
	LessThan1,
	always0,
	always01,
	ccifiwait_0,
	nRST,
	devpor,
	devclrn,
	devoe);
input 	prifdmemren;
input 	prifdmemwen;
input 	LessThan1;
input 	always0;
output 	always01;
output 	ccifiwait_0;
input 	nRST;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X55_Y30_N28
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// always01 = (prifdmemren) # (prifdmemwen)

	.dataa(gnd),
	.datab(gnd),
	.datac(prifdmemren),
	.datad(prifdmemwen),
	.cin(gnd),
	.combout(always01),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'hFFF0;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X55_Y30_N4
cycloneive_lcell_comb \ccif.iwait[0]~0 (
// Equation(s):
// ccifiwait_0 = (always01) # ((\nRST~input_o  & ((!always0) # (!LessThan1))))

	.dataa(nRST),
	.datab(LessThan1),
	.datac(always0),
	.datad(always01),
	.cin(gnd),
	.combout(ccifiwait_0),
	.cout());
// synopsys translate_off
defparam \ccif.iwait[0]~0 .lut_mask = 16'hFF2A;
defparam \ccif.iwait[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module ram (
	is_in_use_reg,
	LessThan1,
	\ramif.ramaddr ,
	ramaddr,
	ramaddr1,
	ramaddr2,
	ramaddr3,
	ramaddr4,
	ramaddr5,
	ramaddr6,
	ramaddr7,
	ramaddr8,
	ramaddr9,
	ramaddr10,
	ramaddr11,
	ramaddr12,
	ramaddr13,
	ramaddr14,
	\ramif.ramWEN ,
	\ramif.ramREN ,
	ramaddr15,
	ramaddr16,
	always0,
	always1,
	ramiframload_0,
	ramiframload_1,
	ramiframload_2,
	ramiframload_3,
	ramiframload_4,
	ramiframload_5,
	ramiframload_6,
	ramiframload_7,
	ramiframload_8,
	ramiframload_9,
	ramiframload_10,
	ramiframload_11,
	ramiframload_12,
	ramiframload_13,
	ramiframload_14,
	ramiframload_15,
	ramiframload_16,
	ramiframload_17,
	ramiframload_18,
	ramiframload_19,
	ramiframload_20,
	ramiframload_21,
	ramiframload_22,
	ramiframload_23,
	ramiframload_24,
	ramiframload_25,
	ramiframload_26,
	ramiframload_27,
	ramiframload_28,
	ramiframload_29,
	ramiframload_30,
	ramiframload_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	ramstore,
	ramstore1,
	ramstore2,
	ramstore3,
	ramstore4,
	ramstore5,
	ramstore6,
	ramstore7,
	ramstore8,
	ramstore9,
	ramstore10,
	ramstore11,
	ramstore12,
	ramstore13,
	ramstore14,
	ramstore15,
	ramstore16,
	ramstore17,
	ramstore18,
	ramstore19,
	ramstore20,
	ramstore21,
	ramstore22,
	ramstore23,
	ramstore24,
	ramstore25,
	ramstore26,
	ramstore27,
	ramstore28,
	ramstore29,
	ramstore30,
	ramstore31,
	ramaddr17,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	nRST,
	altera_internal_jtag1,
	nRST1,
	CLK,
	devpor,
	devclrn,
	devoe);
output 	is_in_use_reg;
output 	LessThan1;
input 	[31:0] \ramif.ramaddr ;
input 	ramaddr;
input 	ramaddr1;
input 	ramaddr2;
input 	ramaddr3;
input 	ramaddr4;
input 	ramaddr5;
input 	ramaddr6;
input 	ramaddr7;
input 	ramaddr8;
input 	ramaddr9;
input 	ramaddr10;
input 	ramaddr11;
input 	ramaddr12;
input 	ramaddr13;
input 	ramaddr14;
input 	\ramif.ramWEN ;
input 	\ramif.ramREN ;
input 	ramaddr15;
input 	ramaddr16;
output 	always0;
output 	always1;
output 	ramiframload_0;
output 	ramiframload_1;
output 	ramiframload_2;
output 	ramiframload_3;
output 	ramiframload_4;
output 	ramiframload_5;
output 	ramiframload_6;
output 	ramiframload_7;
output 	ramiframload_8;
output 	ramiframload_9;
output 	ramiframload_10;
output 	ramiframload_11;
output 	ramiframload_12;
output 	ramiframload_13;
output 	ramiframload_14;
output 	ramiframload_15;
output 	ramiframload_16;
output 	ramiframload_17;
output 	ramiframload_18;
output 	ramiframload_19;
output 	ramiframload_20;
output 	ramiframload_21;
output 	ramiframload_22;
output 	ramiframload_23;
output 	ramiframload_24;
output 	ramiframload_25;
output 	ramiframload_26;
output 	ramiframload_27;
output 	ramiframload_28;
output 	ramiframload_29;
output 	ramiframload_30;
output 	ramiframload_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	ramstore;
input 	ramstore1;
input 	ramstore2;
input 	ramstore3;
input 	ramstore4;
input 	ramstore5;
input 	ramstore6;
input 	ramstore7;
input 	ramstore8;
input 	ramstore9;
input 	ramstore10;
input 	ramstore11;
input 	ramstore12;
input 	ramstore13;
input 	ramstore14;
input 	ramstore15;
input 	ramstore16;
input 	ramstore17;
input 	ramstore18;
input 	ramstore19;
input 	ramstore20;
input 	ramstore21;
input 	ramstore22;
input 	ramstore23;
input 	ramstore24;
input 	ramstore25;
input 	ramstore26;
input 	ramstore27;
input 	ramstore28;
input 	ramstore29;
input 	ramstore30;
input 	ramstore31;
input 	ramaddr17;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	nRST;
input 	altera_internal_jtag1;
input 	nRST1;
input 	CLK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ;
wire \altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ;
wire \always0~1_combout ;
wire \always0~10_combout ;
wire \always0~17_combout ;
wire \always0~22_combout ;
wire \always0~2_combout ;
wire \addr[0]~feeder_combout ;
wire \always0~0_combout ;
wire \always0~3_combout ;
wire \always0~4_combout ;
wire \always0~11_combout ;
wire \always0~13_combout ;
wire \always0~12_combout ;
wire \always0~14_combout ;
wire \always0~15_combout ;
wire \always0~18_combout ;
wire \addr[18]~feeder_combout ;
wire \always0~16_combout ;
wire \always0~19_combout ;
wire \always0~20_combout ;
wire \always0~23_combout ;
wire \count[0]~3_combout ;
wire \count[1]~2_combout ;
wire \Add0~1_combout ;
wire \count[2]~1_combout ;
wire \Add0~0_combout ;
wire \count[3]~0_combout ;
wire \always0~5_combout ;
wire \always0~7_combout ;
wire \always0~8_combout ;
wire \always0~6_combout ;
wire \always0~9_combout ;
wire [1:0] en;
wire [3:0] count;
wire [31:0] addr;
wire [0:0] \altsyncram_component|auto_generated|altsyncram1|address_reg_a ;


altsyncram_1 altsyncram_component(
	.ram_block3a32(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.ram_block3a0(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.ram_block3a33(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.ram_block3a1(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.ram_block3a34(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.ram_block3a2(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.ram_block3a35(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.ram_block3a3(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.ram_block3a36(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.ram_block3a4(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.ram_block3a37(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.ram_block3a5(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.ram_block3a38(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.ram_block3a6(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.ram_block3a39(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.ram_block3a7(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.ram_block3a40(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.ram_block3a8(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.ram_block3a41(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.ram_block3a9(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.ram_block3a42(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.ram_block3a10(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.ram_block3a43(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.ram_block3a11(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.ram_block3a44(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.ram_block3a12(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.ram_block3a45(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.ram_block3a13(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.ram_block3a46(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.ram_block3a14(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.ram_block3a47(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.ram_block3a15(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.ram_block3a48(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.ram_block3a16(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.ram_block3a49(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.ram_block3a17(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.ram_block3a50(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.ram_block3a18(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.ram_block3a51(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.ram_block3a19(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.ram_block3a52(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.ram_block3a20(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.ram_block3a53(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.ram_block3a21(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.ram_block3a54(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.ram_block3a22(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.ram_block3a55(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.ram_block3a23(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.ram_block3a56(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.ram_block3a24(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.ram_block3a57(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.ram_block3a25(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.ram_block3a58(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.ram_block3a26(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.ram_block3a59(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.ram_block3a27(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.ram_block3a60(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.ram_block3a28(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.ram_block3a61(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.ram_block3a29(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.ram_block3a62(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.ram_block3a30(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.ram_block3a63(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.ram_block3a31(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.address_a({gnd,ramaddr14,ramaddr11,ramaddr12,ramaddr9,ramaddr10,ramaddr7,ramaddr8,ramaddr5,ramaddr6,ramaddr3,ramaddr4,ramaddr1,ramaddr2}),
	.ramaddr(ramaddr13),
	.ramWEN(\ramif.ramWEN ),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({ramstore31,ramstore30,ramstore29,ramstore28,ramstore27,ramstore26,ramstore25,ramstore24,ramstore23,ramstore22,ramstore21,ramstore20,ramstore19,ramstore18,ramstore17,ramstore16,ramstore15,ramstore14,ramstore13,ramstore12,ramstore11,ramstore10,ramstore9,ramstore8,ramstore7,ramstore6,
ramstore5,ramstore4,ramstore3,ramstore2,ramstore1,ramstore}),
	.ramaddr1(ramaddr17),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(CLK),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: FF_X60_Y29_N17
dffeas \addr[2] (
	.clk(CLK),
	.d(ramaddr2),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[2]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[2] .is_wysiwyg = "true";
defparam \addr[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X60_Y29_N11
dffeas \addr[3] (
	.clk(CLK),
	.d(ramaddr1),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[3]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[3] .is_wysiwyg = "true";
defparam \addr[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N4
cycloneive_lcell_comb \always0~1 (
// Equation(s):
// \always0~1_combout  = (\ramaddr~5_combout  & (addr[3] & (addr[2] $ (!\ramaddr~7_combout )))) # (!\ramaddr~5_combout  & (!addr[3] & (addr[2] $ (!\ramaddr~7_combout ))))

	.dataa(ramaddr1),
	.datab(addr[3]),
	.datac(addr[2]),
	.datad(ramaddr2),
	.cin(gnd),
	.combout(\always0~1_combout ),
	.cout());
// synopsys translate_off
defparam \always0~1 .lut_mask = 16'h9009;
defparam \always0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y28_N7
dffeas \addr[5] (
	.clk(CLK),
	.d(ramaddr3),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[5]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[5] .is_wysiwyg = "true";
defparam \addr[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X54_Y29_N17
dffeas \addr[6] (
	.clk(CLK),
	.d(ramaddr6),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[6]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[6] .is_wysiwyg = "true";
defparam \addr[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y25_N3
dffeas \addr[10] (
	.clk(CLK),
	.d(ramaddr10),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[10]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[10] .is_wysiwyg = "true";
defparam \addr[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N5
dffeas \addr[13] (
	.clk(CLK),
	.d(ramaddr11),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[13]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[13] .is_wysiwyg = "true";
defparam \addr[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y26_N3
dffeas \addr[14] (
	.clk(CLK),
	.d(ramaddr14),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[14]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[14] .is_wysiwyg = "true";
defparam \addr[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N13
dffeas \addr[22] (
	.clk(CLK),
	.d(\ramif.ramaddr [22]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[22]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[22] .is_wysiwyg = "true";
defparam \addr[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y30_N7
dffeas \addr[23] (
	.clk(CLK),
	.d(\ramif.ramaddr [23]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[23]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[23] .is_wysiwyg = "true";
defparam \addr[23] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y30_N20
cycloneive_lcell_comb \always0~10 (
// Equation(s):
// \always0~10_combout  = (\ramaddr~35_combout  & (addr[22] & (addr[23] $ (!\ramaddr~33_combout )))) # (!\ramaddr~35_combout  & (!addr[22] & (addr[23] $ (!\ramaddr~33_combout ))))

	.dataa(\ramif.ramaddr [22]),
	.datab(addr[23]),
	.datac(addr[22]),
	.datad(\ramif.ramaddr [23]),
	.cin(gnd),
	.combout(\always0~10_combout ),
	.cout());
// synopsys translate_off
defparam \always0~10 .lut_mask = 16'h8421;
defparam \always0~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y29_N7
dffeas \addr[29] (
	.clk(CLK),
	.d(\ramif.ramaddr [29]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[29]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[29] .is_wysiwyg = "true";
defparam \addr[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y29_N1
dffeas \addr[31] (
	.clk(CLK),
	.d(\ramif.ramaddr [31]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[31]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[31] .is_wysiwyg = "true";
defparam \addr[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y31_N23
dffeas \addr[20] (
	.clk(CLK),
	.d(\ramif.ramaddr [20]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[20]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[20] .is_wysiwyg = "true";
defparam \addr[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X61_Y29_N17
dffeas \addr[17] (
	.clk(CLK),
	.d(\ramif.ramaddr [17]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[17]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[17] .is_wysiwyg = "true";
defparam \addr[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X55_Y29_N29
dffeas \addr[19] (
	.clk(CLK),
	.d(\ramif.ramaddr [19]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[19]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[19] .is_wysiwyg = "true";
defparam \addr[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y29_N19
dffeas \addr[24] (
	.clk(CLK),
	.d(gnd),
	.asdata(ramaddr16),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[24]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[24] .is_wysiwyg = "true";
defparam \addr[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X58_Y29_N17
dffeas \addr[25] (
	.clk(CLK),
	.d(\ramif.ramaddr [25]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[25]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[25] .is_wysiwyg = "true";
defparam \addr[25] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N12
cycloneive_lcell_comb \always0~17 (
// Equation(s):
// \always0~17_combout  = (addr[25] & (\ramaddr~57_combout  & (addr[24] $ (!\ramaddr~59_combout )))) # (!addr[25] & (!\ramaddr~57_combout  & (addr[24] $ (!\ramaddr~59_combout ))))

	.dataa(addr[25]),
	.datab(addr[24]),
	.datac(\ramif.ramaddr [25]),
	.datad(ramaddr16),
	.cin(gnd),
	.combout(\always0~17_combout ),
	.cout());
// synopsys translate_off
defparam \always0~17 .lut_mask = 16'h8421;
defparam \always0~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N14
cycloneive_lcell_comb \LessThan1~0 (
// Equation(s):
// LessThan1 = (count[2]) # ((count[3]) # (count[1]))

	.dataa(count[2]),
	.datab(count[3]),
	.datac(count[1]),
	.datad(gnd),
	.cin(gnd),
	.combout(LessThan1),
	.cout());
// synopsys translate_off
defparam \LessThan1~0 .lut_mask = 16'hFEFE;
defparam \LessThan1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N16
cycloneive_lcell_comb \always0~21 (
// Equation(s):
// always0 = (\always0~4_combout  & (\always0~9_combout  & \always0~20_combout ))

	.dataa(\always0~4_combout ),
	.datab(\always0~9_combout ),
	.datac(gnd),
	.datad(\always0~20_combout ),
	.cin(gnd),
	.combout(always0),
	.cout());
// synopsys translate_off
defparam \always0~21 .lut_mask = 16'h8800;
defparam \always0~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N18
cycloneive_lcell_comb \always1~0 (
// Equation(s):
// always1 = ((LessThan1 & always0)) # (!\nRST~input_o )

	.dataa(nRST),
	.datab(LessThan1),
	.datac(gnd),
	.datad(always0),
	.cin(gnd),
	.combout(always1),
	.cout());
// synopsys translate_off
defparam \always1~0 .lut_mask = 16'hDD55;
defparam \always1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y28_N24
cycloneive_lcell_comb \ramif.ramload[0]~0 (
// Equation(s):
// ramiframload_0 = ((address_reg_a_0 & (ram_block3a321)) # (!address_reg_a_0 & ((ram_block3a01)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a32~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a0~portadataout ),
	.datad(always1),
	.cin(gnd),
	.combout(ramiframload_0),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[0]~0 .lut_mask = 16'hD8FF;
defparam \ramif.ramload[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N10
cycloneive_lcell_comb \ramif.ramload[1]~1 (
// Equation(s):
// ramiframload_1 = (always1 & ((address_reg_a_0 & (ram_block3a331)) # (!address_reg_a_0 & ((ram_block3a110)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a33~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a1~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_1),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[1]~1 .lut_mask = 16'hA0C0;
defparam \ramif.ramload[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N6
cycloneive_lcell_comb \ramif.ramload[2]~2 (
// Equation(s):
// ramiframload_2 = (always1 & ((address_reg_a_0 & (ram_block3a341)) # (!address_reg_a_0 & ((ram_block3a210)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a34~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a2~portadataout ),
	.cin(gnd),
	.combout(ramiframload_2),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[2]~2 .lut_mask = 16'hC480;
defparam \ramif.ramload[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N0
cycloneive_lcell_comb \ramif.ramload[3]~3 (
// Equation(s):
// ramiframload_3 = (always1 & ((address_reg_a_0 & ((ram_block3a351))) # (!address_reg_a_0 & (ram_block3a310))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a3~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a35~portadataout ),
	.cin(gnd),
	.combout(ramiframload_3),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[3]~3 .lut_mask = 16'hC808;
defparam \ramif.ramload[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y27_N22
cycloneive_lcell_comb \ramif.ramload[4]~4 (
// Equation(s):
// ramiframload_4 = ((address_reg_a_0 & ((ram_block3a361))) # (!address_reg_a_0 & (ram_block3a410))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a4~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a36~portadataout ),
	.cin(gnd),
	.combout(ramiframload_4),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[4]~4 .lut_mask = 16'hEF4F;
defparam \ramif.ramload[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N6
cycloneive_lcell_comb \ramif.ramload[5]~5 (
// Equation(s):
// ramiframload_5 = (always1 & ((address_reg_a_0 & ((ram_block3a371))) # (!address_reg_a_0 & (ram_block3a510))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a5~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a37~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_5),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[5]~5 .lut_mask = 16'hC088;
defparam \ramif.ramload[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N24
cycloneive_lcell_comb \ramif.ramload[6]~6 (
// Equation(s):
// ramiframload_6 = ((address_reg_a_0 & ((ram_block3a381))) # (!address_reg_a_0 & (ram_block3a64))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a6~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a38~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_6),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[6]~6 .lut_mask = 16'hCFAF;
defparam \ramif.ramload[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N20
cycloneive_lcell_comb \ramif.ramload[7]~7 (
// Equation(s):
// ramiframload_7 = ((address_reg_a_0 & ((ram_block3a391))) # (!address_reg_a_0 & (ram_block3a71))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a7~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a39~portadataout ),
	.cin(gnd),
	.combout(ramiframload_7),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[7]~7 .lut_mask = 16'hEF2F;
defparam \ramif.ramload[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N26
cycloneive_lcell_comb \ramif.ramload[8]~8 (
// Equation(s):
// ramiframload_8 = (always1 & ((address_reg_a_0 & ((ram_block3a401))) # (!address_reg_a_0 & (ram_block3a81))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a8~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a40~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_8),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[8]~8 .lut_mask = 16'hC0A0;
defparam \ramif.ramload[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N26
cycloneive_lcell_comb \ramif.ramload[9]~9 (
// Equation(s):
// ramiframload_9 = ((address_reg_a_0 & ((ram_block3a412))) # (!address_reg_a_0 & (ram_block3a91))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a9~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a41~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_9),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[9]~9 .lut_mask = 16'hCFAF;
defparam \ramif.ramload[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N24
cycloneive_lcell_comb \ramif.ramload[10]~10 (
// Equation(s):
// ramiframload_10 = (always1 & ((address_reg_a_0 & ((ram_block3a421))) # (!address_reg_a_0 & (ram_block3a101))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a10~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a42~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_10),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[10]~10 .lut_mask = 16'hC0A0;
defparam \ramif.ramload[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N10
cycloneive_lcell_comb \ramif.ramload[11]~11 (
// Equation(s):
// ramiframload_11 = ((address_reg_a_0 & (ram_block3a431)) # (!address_reg_a_0 & ((ram_block3a112)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a43~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a11~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_11),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[11]~11 .lut_mask = 16'hBBF3;
defparam \ramif.ramload[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N16
cycloneive_lcell_comb \ramif.ramload[12]~12 (
// Equation(s):
// ramiframload_12 = ((address_reg_a_0 & (ram_block3a441)) # (!address_reg_a_0 & ((ram_block3a121)))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a44~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a12~portadataout ),
	.cin(gnd),
	.combout(ramiframload_12),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[12]~12 .lut_mask = 16'hBF8F;
defparam \ramif.ramload[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N22
cycloneive_lcell_comb \ramif.ramload[13]~13 (
// Equation(s):
// ramiframload_13 = ((address_reg_a_0 & ((ram_block3a451))) # (!address_reg_a_0 & (ram_block3a131))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a13~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a45~portadataout ),
	.cin(gnd),
	.combout(ramiframload_13),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[13]~13 .lut_mask = 16'hFD75;
defparam \ramif.ramload[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N12
cycloneive_lcell_comb \ramif.ramload[14]~14 (
// Equation(s):
// ramiframload_14 = (always1 & ((address_reg_a_0 & ((ram_block3a461))) # (!address_reg_a_0 & (ram_block3a141))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a14~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a46~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_14),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[14]~14 .lut_mask = 16'hC088;
defparam \ramif.ramload[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N12
cycloneive_lcell_comb \ramif.ramload[15]~15 (
// Equation(s):
// ramiframload_15 = ((address_reg_a_0 & ((ram_block3a471))) # (!address_reg_a_0 & (ram_block3a151))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a15~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a47~portadataout ),
	.cin(gnd),
	.combout(ramiframload_15),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[15]~15 .lut_mask = 16'hFD75;
defparam \ramif.ramload[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N6
cycloneive_lcell_comb \ramif.ramload[16]~16 (
// Equation(s):
// ramiframload_16 = ((address_reg_a_0 & (ram_block3a481)) # (!address_reg_a_0 & ((ram_block3a161)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a48~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a16~portadataout ),
	.cin(gnd),
	.combout(ramiframload_16),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[16]~16 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N20
cycloneive_lcell_comb \ramif.ramload[17]~17 (
// Equation(s):
// ramiframload_17 = (always1 & ((address_reg_a_0 & ((ram_block3a491))) # (!address_reg_a_0 & (ram_block3a171))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a17~portadataout ),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a49~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_17),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[17]~17 .lut_mask = 16'hA088;
defparam \ramif.ramload[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y30_N10
cycloneive_lcell_comb \ramif.ramload[18]~18 (
// Equation(s):
// ramiframload_18 = (always1 & ((address_reg_a_0 & ((ram_block3a501))) # (!address_reg_a_0 & (ram_block3a181))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a18~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a50~portadataout ),
	.cin(gnd),
	.combout(ramiframload_18),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[18]~18 .lut_mask = 16'hE020;
defparam \ramif.ramload[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N30
cycloneive_lcell_comb \ramif.ramload[19]~19 (
// Equation(s):
// ramiframload_19 = (always1 & ((address_reg_a_0 & ((ram_block3a512))) # (!address_reg_a_0 & (ram_block3a191))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a19~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a51~portadataout ),
	.cin(gnd),
	.combout(ramiframload_19),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[19]~19 .lut_mask = 16'hE020;
defparam \ramif.ramload[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N10
cycloneive_lcell_comb \ramif.ramload[20]~20 (
// Equation(s):
// ramiframload_20 = ((address_reg_a_0 & ((ram_block3a521))) # (!address_reg_a_0 & (ram_block3a201))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a20~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a52~portadataout ),
	.cin(gnd),
	.combout(ramiframload_20),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[20]~20 .lut_mask = 16'hFD75;
defparam \ramif.ramload[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N8
cycloneive_lcell_comb \ramif.ramload[21]~21 (
// Equation(s):
// ramiframload_21 = (always1 & ((address_reg_a_0 & (ram_block3a531)) # (!address_reg_a_0 & ((ram_block3a212)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a53~portadataout ),
	.datab(always1),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a21~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_21),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[21]~21 .lut_mask = 16'h88C0;
defparam \ramif.ramload[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N10
cycloneive_lcell_comb \ramif.ramload[22]~22 (
// Equation(s):
// ramiframload_22 = ((address_reg_a_0 & ((ram_block3a541))) # (!address_reg_a_0 & (ram_block3a221))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a22~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a54~portadataout ),
	.cin(gnd),
	.combout(ramiframload_22),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[22]~22 .lut_mask = 16'hFD75;
defparam \ramif.ramload[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N24
cycloneive_lcell_comb \ramif.ramload[23]~23 (
// Equation(s):
// ramiframload_23 = ((address_reg_a_0 & (ram_block3a551)) # (!address_reg_a_0 & ((ram_block3a231)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a55~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a23~portadataout ),
	.cin(gnd),
	.combout(ramiframload_23),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[23]~23 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y32_N30
cycloneive_lcell_comb \ramif.ramload[24]~24 (
// Equation(s):
// ramiframload_24 = (always1 & ((address_reg_a_0 & (ram_block3a561)) # (!address_reg_a_0 & ((ram_block3a241)))))

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a56~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a24~portadataout ),
	.cin(gnd),
	.combout(ramiframload_24),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[24]~24 .lut_mask = 16'hB080;
defparam \ramif.ramload[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y28_N0
cycloneive_lcell_comb \ramif.ramload[25]~25 (
// Equation(s):
// ramiframload_25 = ((address_reg_a_0 & ((ram_block3a571))) # (!address_reg_a_0 & (ram_block3a251))) # (!always1)

	.dataa(\altsyncram_component|auto_generated|altsyncram1|ram_block3a25~portadataout ),
	.datab(\altsyncram_component|auto_generated|altsyncram1|ram_block3a57~portadataout ),
	.datac(always1),
	.datad(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.cin(gnd),
	.combout(ramiframload_25),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[25]~25 .lut_mask = 16'hCFAF;
defparam \ramif.ramload[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N12
cycloneive_lcell_comb \ramif.ramload[26]~26 (
// Equation(s):
// ramiframload_26 = (always1 & ((address_reg_a_0 & ((ram_block3a581))) # (!address_reg_a_0 & (ram_block3a261))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a26~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a58~portadataout ),
	.cin(gnd),
	.combout(ramiframload_26),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[26]~26 .lut_mask = 16'hA820;
defparam \ramif.ramload[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N30
cycloneive_lcell_comb \ramif.ramload[27]~27 (
// Equation(s):
// ramiframload_27 = ((address_reg_a_0 & ((ram_block3a591))) # (!address_reg_a_0 & (ram_block3a271))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a27~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a59~portadataout ),
	.cin(gnd),
	.combout(ramiframload_27),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[27]~27 .lut_mask = 16'hFD75;
defparam \ramif.ramload[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N0
cycloneive_lcell_comb \ramif.ramload[28]~28 (
// Equation(s):
// ramiframload_28 = ((address_reg_a_0 & (ram_block3a601)) # (!address_reg_a_0 & ((ram_block3a281)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a60~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a28~portadataout ),
	.cin(gnd),
	.combout(ramiframload_28),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[28]~28 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N26
cycloneive_lcell_comb \ramif.ramload[29]~29 (
// Equation(s):
// ramiframload_29 = ((address_reg_a_0 & (ram_block3a611)) # (!address_reg_a_0 & ((ram_block3a291)))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a61~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a29~portadataout ),
	.cin(gnd),
	.combout(ramiframload_29),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[29]~29 .lut_mask = 16'hF7D5;
defparam \ramif.ramload[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N8
cycloneive_lcell_comb \ramif.ramload[30]~30 (
// Equation(s):
// ramiframload_30 = (always1 & ((address_reg_a_0 & (ram_block3a621)) # (!address_reg_a_0 & ((ram_block3a301)))))

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a62~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a30~portadataout ),
	.cin(gnd),
	.combout(ramiframload_30),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[30]~30 .lut_mask = 16'hA280;
defparam \ramif.ramload[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X53_Y31_N18
cycloneive_lcell_comb \ramif.ramload[31]~31 (
// Equation(s):
// ramiframload_31 = ((address_reg_a_0 & ((ram_block3a631))) # (!address_reg_a_0 & (ram_block3a312))) # (!always1)

	.dataa(always1),
	.datab(\altsyncram_component|auto_generated|altsyncram1|address_reg_a [0]),
	.datac(\altsyncram_component|auto_generated|altsyncram1|ram_block3a31~portadataout ),
	.datad(\altsyncram_component|auto_generated|altsyncram1|ram_block3a63~portadataout ),
	.cin(gnd),
	.combout(ramiframload_31),
	.cout());
// synopsys translate_off
defparam \ramif.ramload[31]~31 .lut_mask = 16'hFD75;
defparam \ramif.ramload[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y29_N23
dffeas \en[0] (
	.clk(CLK),
	.d(\ramif.ramWEN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[0]),
	.prn(vcc));
// synopsys translate_off
defparam \en[0] .is_wysiwyg = "true";
defparam \en[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X62_Y29_N5
dffeas \en[1] (
	.clk(CLK),
	.d(\ramif.ramREN ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(en[1]),
	.prn(vcc));
// synopsys translate_off
defparam \en[1] .is_wysiwyg = "true";
defparam \en[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N8
cycloneive_lcell_comb \always0~22 (
// Equation(s):
// \always0~22_combout  = (\ramWEN~0_combout  & ((\ramREN~0_combout  $ (en[1])) # (!en[0]))) # (!\ramWEN~0_combout  & ((en[0]) # (\ramREN~0_combout  $ (en[1]))))

	.dataa(\ramif.ramWEN ),
	.datab(en[0]),
	.datac(\ramif.ramREN ),
	.datad(en[1]),
	.cin(gnd),
	.combout(\always0~22_combout ),
	.cout());
// synopsys translate_off
defparam \always0~22 .lut_mask = 16'h6FF6;
defparam \always0~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y28_N5
dffeas \addr[4] (
	.clk(CLK),
	.d(ramaddr4),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[4]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[4] .is_wysiwyg = "true";
defparam \addr[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y28_N0
cycloneive_lcell_comb \always0~2 (
// Equation(s):
// \always0~2_combout  = (addr[5] & (\ramaddr~9_combout  & (addr[4] $ (!\ramaddr~11_combout )))) # (!addr[5] & (!\ramaddr~9_combout  & (addr[4] $ (!\ramaddr~11_combout ))))

	.dataa(addr[5]),
	.datab(addr[4]),
	.datac(ramaddr4),
	.datad(ramaddr3),
	.cin(gnd),
	.combout(\always0~2_combout ),
	.cout());
// synopsys translate_off
defparam \always0~2 .lut_mask = 16'h8241;
defparam \always0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y29_N3
dffeas \addr[1] (
	.clk(CLK),
	.d(\ramif.ramaddr [1]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[1]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[1] .is_wysiwyg = "true";
defparam \addr[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N20
cycloneive_lcell_comb \addr[0]~feeder (
// Equation(s):
// \addr[0]~feeder_combout  = \ramaddr~3_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ramaddr),
	.cin(gnd),
	.combout(\addr[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[0]~feeder .lut_mask = 16'hFF00;
defparam \addr[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y29_N21
dffeas \addr[0] (
	.clk(CLK),
	.d(\addr[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[0]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[0] .is_wysiwyg = "true";
defparam \addr[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y29_N14
cycloneive_lcell_comb \always0~0 (
// Equation(s):
// \always0~0_combout  = (\ramaddr~3_combout  & (addr[0] & (addr[1] $ (!\ramaddr~1_combout )))) # (!\ramaddr~3_combout  & (!addr[0] & (addr[1] $ (!\ramaddr~1_combout ))))

	.dataa(ramaddr),
	.datab(addr[1]),
	.datac(addr[0]),
	.datad(\ramif.ramaddr [1]),
	.cin(gnd),
	.combout(\always0~0_combout ),
	.cout());
// synopsys translate_off
defparam \always0~0 .lut_mask = 16'h8421;
defparam \always0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X54_Y29_N23
dffeas \addr[7] (
	.clk(CLK),
	.d(ramaddr5),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[7]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[7] .is_wysiwyg = "true";
defparam \addr[7] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X54_Y29_N12
cycloneive_lcell_comb \always0~3 (
// Equation(s):
// \always0~3_combout  = (addr[6] & (\ramaddr~15_combout  & (addr[7] $ (!\ramaddr~13_combout )))) # (!addr[6] & (!\ramaddr~15_combout  & (addr[7] $ (!\ramaddr~13_combout ))))

	.dataa(addr[6]),
	.datab(addr[7]),
	.datac(ramaddr5),
	.datad(ramaddr6),
	.cin(gnd),
	.combout(\always0~3_combout ),
	.cout());
// synopsys translate_off
defparam \always0~3 .lut_mask = 16'h8241;
defparam \always0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N30
cycloneive_lcell_comb \always0~4 (
// Equation(s):
// \always0~4_combout  = (\always0~1_combout  & (\always0~2_combout  & (\always0~0_combout  & \always0~3_combout )))

	.dataa(\always0~1_combout ),
	.datab(\always0~2_combout ),
	.datac(\always0~0_combout ),
	.datad(\always0~3_combout ),
	.cin(gnd),
	.combout(\always0~4_combout ),
	.cout());
// synopsys translate_off
defparam \always0~4 .lut_mask = 16'h8000;
defparam \always0~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X62_Y29_N11
dffeas \addr[21] (
	.clk(CLK),
	.d(\ramif.ramaddr [21]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[21]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[21] .is_wysiwyg = "true";
defparam \addr[21] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X62_Y29_N2
cycloneive_lcell_comb \always0~11 (
// Equation(s):
// \always0~11_combout  = (\ramWEN~0_combout  & (!\ramREN~0_combout  & (addr[21] $ (!\ramaddr~37_combout )))) # (!\ramWEN~0_combout  & (addr[21] $ (((!\ramaddr~37_combout )))))

	.dataa(\ramif.ramWEN ),
	.datab(addr[21]),
	.datac(\ramif.ramREN ),
	.datad(\ramif.ramaddr [21]),
	.cin(gnd),
	.combout(\always0~11_combout ),
	.cout());
// synopsys translate_off
defparam \always0~11 .lut_mask = 16'h4C13;
defparam \always0~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y29_N23
dffeas \addr[30] (
	.clk(CLK),
	.d(\ramif.ramaddr [30]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[30]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[30] .is_wysiwyg = "true";
defparam \addr[30] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N26
cycloneive_lcell_comb \always0~13 (
// Equation(s):
// \always0~13_combout  = (addr[31] & (\ramaddr~43_combout  & (addr[30] $ (!\ramaddr~45_combout )))) # (!addr[31] & (!\ramaddr~43_combout  & (addr[30] $ (!\ramaddr~45_combout ))))

	.dataa(addr[31]),
	.datab(addr[30]),
	.datac(\ramif.ramaddr [30]),
	.datad(\ramif.ramaddr [31]),
	.cin(gnd),
	.combout(\always0~13_combout ),
	.cout());
// synopsys translate_off
defparam \always0~13 .lut_mask = 16'h8241;
defparam \always0~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X58_Y29_N5
dffeas \addr[28] (
	.clk(CLK),
	.d(\ramif.ramaddr [28]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[28]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[28] .is_wysiwyg = "true";
defparam \addr[28] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X58_Y29_N8
cycloneive_lcell_comb \always0~12 (
// Equation(s):
// \always0~12_combout  = (addr[29] & (\ramaddr~39_combout  & (addr[28] $ (!\ramaddr~41_combout )))) # (!addr[29] & (!\ramaddr~39_combout  & (addr[28] $ (!\ramaddr~41_combout ))))

	.dataa(addr[29]),
	.datab(addr[28]),
	.datac(\ramif.ramaddr [28]),
	.datad(\ramif.ramaddr [29]),
	.cin(gnd),
	.combout(\always0~12_combout ),
	.cout());
// synopsys translate_off
defparam \always0~12 .lut_mask = 16'h8241;
defparam \always0~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N8
cycloneive_lcell_comb \always0~14 (
// Equation(s):
// \always0~14_combout  = (\always0~13_combout  & (\always0~12_combout  & (addr[20] $ (!\ramaddr~47_combout ))))

	.dataa(addr[20]),
	.datab(\ramif.ramaddr [20]),
	.datac(\always0~13_combout ),
	.datad(\always0~12_combout ),
	.cin(gnd),
	.combout(\always0~14_combout ),
	.cout());
// synopsys translate_off
defparam \always0~14 .lut_mask = 16'h9000;
defparam \always0~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X61_Y29_N31
dffeas \addr[16] (
	.clk(CLK),
	.d(\ramif.ramaddr [16]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[16]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[16] .is_wysiwyg = "true";
defparam \addr[16] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X61_Y29_N2
cycloneive_lcell_comb \always0~15 (
// Equation(s):
// \always0~15_combout  = (addr[17] & (\ramaddr~49_combout  & (addr[16] $ (!\ramaddr~51_combout )))) # (!addr[17] & (!\ramaddr~49_combout  & (addr[16] $ (!\ramaddr~51_combout ))))

	.dataa(addr[17]),
	.datab(addr[16]),
	.datac(\ramif.ramaddr [16]),
	.datad(\ramif.ramaddr [17]),
	.cin(gnd),
	.combout(\always0~15_combout ),
	.cout());
// synopsys translate_off
defparam \always0~15 .lut_mask = 16'h8241;
defparam \always0~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y29_N21
dffeas \addr[27] (
	.clk(CLK),
	.d(\ramif.ramaddr [27]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[27]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[27] .is_wysiwyg = "true";
defparam \addr[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X59_Y29_N7
dffeas \addr[26] (
	.clk(CLK),
	.d(\ramif.ramaddr [26]),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[26]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[26] .is_wysiwyg = "true";
defparam \addr[26] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N26
cycloneive_lcell_comb \always0~18 (
// Equation(s):
// \always0~18_combout  = (\ramaddr~63_combout  & (addr[26] & (addr[27] $ (!\ramaddr~61_combout )))) # (!\ramaddr~63_combout  & (!addr[26] & (addr[27] $ (!\ramaddr~61_combout ))))

	.dataa(\ramif.ramaddr [26]),
	.datab(addr[27]),
	.datac(addr[26]),
	.datad(\ramif.ramaddr [27]),
	.cin(gnd),
	.combout(\always0~18_combout ),
	.cout());
// synopsys translate_off
defparam \always0~18 .lut_mask = 16'h8421;
defparam \always0~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N6
cycloneive_lcell_comb \addr[18]~feeder (
// Equation(s):
// \addr[18]~feeder_combout  = \ramaddr~55_combout 

	.dataa(gnd),
	.datab(gnd),
	.datac(ramaddr15),
	.datad(gnd),
	.cin(gnd),
	.combout(\addr[18]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \addr[18]~feeder .lut_mask = 16'hF0F0;
defparam \addr[18]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X56_Y29_N7
dffeas \addr[18] (
	.clk(CLK),
	.d(\addr[18]~feeder_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[18]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[18] .is_wysiwyg = "true";
defparam \addr[18] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X56_Y29_N16
cycloneive_lcell_comb \always0~16 (
// Equation(s):
// \always0~16_combout  = (addr[19] & (\ramaddr~53_combout  & (addr[18] $ (!\ramaddr~55_combout )))) # (!addr[19] & (!\ramaddr~53_combout  & (addr[18] $ (!\ramaddr~55_combout ))))

	.dataa(addr[19]),
	.datab(addr[18]),
	.datac(ramaddr15),
	.datad(\ramif.ramaddr [19]),
	.cin(gnd),
	.combout(\always0~16_combout ),
	.cout());
// synopsys translate_off
defparam \always0~16 .lut_mask = 16'h8241;
defparam \always0~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N28
cycloneive_lcell_comb \always0~19 (
// Equation(s):
// \always0~19_combout  = (\always0~17_combout  & (\always0~15_combout  & (\always0~18_combout  & \always0~16_combout )))

	.dataa(\always0~17_combout ),
	.datab(\always0~15_combout ),
	.datac(\always0~18_combout ),
	.datad(\always0~16_combout ),
	.cin(gnd),
	.combout(\always0~19_combout ),
	.cout());
// synopsys translate_off
defparam \always0~19 .lut_mask = 16'h8000;
defparam \always0~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N2
cycloneive_lcell_comb \always0~20 (
// Equation(s):
// \always0~20_combout  = (\always0~10_combout  & (\always0~11_combout  & (\always0~14_combout  & \always0~19_combout )))

	.dataa(\always0~10_combout ),
	.datab(\always0~11_combout ),
	.datac(\always0~14_combout ),
	.datad(\always0~19_combout ),
	.cin(gnd),
	.combout(\always0~20_combout ),
	.cout());
// synopsys translate_off
defparam \always0~20 .lut_mask = 16'h8000;
defparam \always0~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N14
cycloneive_lcell_comb \always0~23 (
// Equation(s):
// \always0~23_combout  = ((\always0~22_combout ) # ((!\always0~20_combout ) # (!\always0~4_combout ))) # (!\always0~9_combout )

	.dataa(\always0~9_combout ),
	.datab(\always0~22_combout ),
	.datac(\always0~4_combout ),
	.datad(\always0~20_combout ),
	.cin(gnd),
	.combout(\always0~23_combout ),
	.cout());
// synopsys translate_off
defparam \always0~23 .lut_mask = 16'hDFFF;
defparam \always0~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N0
cycloneive_lcell_comb \count[0]~3 (
// Equation(s):
// \count[0]~3_combout  = (!\always0~23_combout  & (count[0] $ (!LessThan1)))

	.dataa(gnd),
	.datab(\always0~23_combout ),
	.datac(count[0]),
	.datad(LessThan1),
	.cin(gnd),
	.combout(\count[0]~3_combout ),
	.cout());
// synopsys translate_off
defparam \count[0]~3 .lut_mask = 16'h3003;
defparam \count[0]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y29_N1
dffeas \count[0] (
	.clk(CLK),
	.d(\count[0]~3_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[0]),
	.prn(vcc));
// synopsys translate_off
defparam \count[0] .is_wysiwyg = "true";
defparam \count[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N4
cycloneive_lcell_comb \count[1]~2 (
// Equation(s):
// \count[1]~2_combout  = (!\always0~23_combout  & (count[1] $ (((!LessThan1 & count[0])))))

	.dataa(LessThan1),
	.datab(count[0]),
	.datac(count[1]),
	.datad(\always0~23_combout ),
	.cin(gnd),
	.combout(\count[1]~2_combout ),
	.cout());
// synopsys translate_off
defparam \count[1]~2 .lut_mask = 16'h00B4;
defparam \count[1]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N5
dffeas \count[1] (
	.clk(CLK),
	.d(\count[1]~2_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[1]),
	.prn(vcc));
// synopsys translate_off
defparam \count[1] .is_wysiwyg = "true";
defparam \count[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N16
cycloneive_lcell_comb \Add0~1 (
// Equation(s):
// \Add0~1_combout  = count[2] $ (((count[1] & count[0])))

	.dataa(count[2]),
	.datab(gnd),
	.datac(count[1]),
	.datad(count[0]),
	.cin(gnd),
	.combout(\Add0~1_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~1 .lut_mask = 16'h5AAA;
defparam \Add0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N22
cycloneive_lcell_comb \count[2]~1 (
// Equation(s):
// \count[2]~1_combout  = (!\always0~23_combout  & ((LessThan1 & ((count[2]))) # (!LessThan1 & (\Add0~1_combout ))))

	.dataa(LessThan1),
	.datab(\Add0~1_combout ),
	.datac(count[2]),
	.datad(\always0~23_combout ),
	.cin(gnd),
	.combout(\count[2]~1_combout ),
	.cout());
// synopsys translate_off
defparam \count[2]~1 .lut_mask = 16'h00E4;
defparam \count[2]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N23
dffeas \count[2] (
	.clk(CLK),
	.d(\count[2]~1_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[2]),
	.prn(vcc));
// synopsys translate_off
defparam \count[2] .is_wysiwyg = "true";
defparam \count[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N18
cycloneive_lcell_comb \Add0~0 (
// Equation(s):
// \Add0~0_combout  = count[3] $ (((count[1] & (count[0] & count[2]))))

	.dataa(count[1]),
	.datab(count[0]),
	.datac(count[2]),
	.datad(count[3]),
	.cin(gnd),
	.combout(\Add0~0_combout ),
	.cout());
// synopsys translate_off
defparam \Add0~0 .lut_mask = 16'h7F80;
defparam \Add0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X60_Y30_N0
cycloneive_lcell_comb \count[3]~0 (
// Equation(s):
// \count[3]~0_combout  = (!\always0~23_combout  & ((LessThan1 & ((count[3]))) # (!LessThan1 & (\Add0~0_combout ))))

	.dataa(LessThan1),
	.datab(\Add0~0_combout ),
	.datac(count[3]),
	.datad(\always0~23_combout ),
	.cin(gnd),
	.combout(\count[3]~0_combout ),
	.cout());
// synopsys translate_off
defparam \count[3]~0 .lut_mask = 16'h00E4;
defparam \count[3]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X60_Y30_N1
dffeas \count[3] (
	.clk(CLK),
	.d(\count[3]~0_combout ),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(count[3]),
	.prn(vcc));
// synopsys translate_off
defparam \count[3] .is_wysiwyg = "true";
defparam \count[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N27
dffeas \addr[9] (
	.clk(CLK),
	.d(ramaddr7),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[9]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[9] .is_wysiwyg = "true";
defparam \addr[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X57_Y29_N1
dffeas \addr[8] (
	.clk(CLK),
	.d(ramaddr8),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[8]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[8] .is_wysiwyg = "true";
defparam \addr[8] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N20
cycloneive_lcell_comb \always0~5 (
// Equation(s):
// \always0~5_combout  = (\ramaddr~17_combout  & (addr[9] & (addr[8] $ (!\ramaddr~19_combout )))) # (!\ramaddr~17_combout  & (!addr[9] & (addr[8] $ (!\ramaddr~19_combout ))))

	.dataa(ramaddr7),
	.datab(addr[9]),
	.datac(addr[8]),
	.datad(ramaddr8),
	.cin(gnd),
	.combout(\always0~5_combout ),
	.cout());
// synopsys translate_off
defparam \always0~5 .lut_mask = 16'h9009;
defparam \always0~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X57_Y29_N7
dffeas \addr[12] (
	.clk(CLK),
	.d(ramaddr12),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[12]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[12] .is_wysiwyg = "true";
defparam \addr[12] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X57_Y29_N14
cycloneive_lcell_comb \always0~7 (
// Equation(s):
// \always0~7_combout  = (addr[13] & (\ramaddr~25_combout  & (addr[12] $ (!\ramaddr~27_combout )))) # (!addr[13] & (!\ramaddr~25_combout  & (addr[12] $ (!\ramaddr~27_combout ))))

	.dataa(addr[13]),
	.datab(ramaddr11),
	.datac(addr[12]),
	.datad(ramaddr12),
	.cin(gnd),
	.combout(\always0~7_combout ),
	.cout());
// synopsys translate_off
defparam \always0~7 .lut_mask = 16'h9009;
defparam \always0~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y29_N5
dffeas \addr[15] (
	.clk(CLK),
	.d(ramaddr17),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[15]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[15] .is_wysiwyg = "true";
defparam \addr[15] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y26_N16
cycloneive_lcell_comb \always0~8 (
// Equation(s):
// \always0~8_combout  = (addr[14] & (\ramaddr~31_combout  & (addr[15] $ (\ramaddr~29_combout )))) # (!addr[14] & (!\ramaddr~31_combout  & (addr[15] $ (\ramaddr~29_combout ))))

	.dataa(addr[14]),
	.datab(addr[15]),
	.datac(ramaddr13),
	.datad(ramaddr14),
	.cin(gnd),
	.combout(\always0~8_combout ),
	.cout());
// synopsys translate_off
defparam \always0~8 .lut_mask = 16'h2814;
defparam \always0~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X59_Y25_N29
dffeas \addr[11] (
	.clk(CLK),
	.d(ramaddr9),
	.asdata(vcc),
	.clrn(nRST1),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\always0~23_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(addr[11]),
	.prn(vcc));
// synopsys translate_off
defparam \addr[11] .is_wysiwyg = "true";
defparam \addr[11] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X59_Y25_N18
cycloneive_lcell_comb \always0~6 (
// Equation(s):
// \always0~6_combout  = (addr[10] & (\ramaddr~23_combout  & (\ramaddr~21_combout  $ (!addr[11])))) # (!addr[10] & (!\ramaddr~23_combout  & (\ramaddr~21_combout  $ (!addr[11]))))

	.dataa(addr[10]),
	.datab(ramaddr9),
	.datac(addr[11]),
	.datad(ramaddr10),
	.cin(gnd),
	.combout(\always0~6_combout ),
	.cout());
// synopsys translate_off
defparam \always0~6 .lut_mask = 16'h8241;
defparam \always0~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N10
cycloneive_lcell_comb \always0~9 (
// Equation(s):
// \always0~9_combout  = (\always0~5_combout  & (\always0~7_combout  & (\always0~8_combout  & \always0~6_combout )))

	.dataa(\always0~5_combout ),
	.datab(\always0~7_combout ),
	.datac(\always0~8_combout ),
	.datad(\always0~6_combout ),
	.cin(gnd),
	.combout(\always0~9_combout ),
	.cout());
// synopsys translate_off
defparam \always0~9 .lut_mask = 16'h8000;
defparam \always0~9 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module altsyncram_1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



altsyncram_99f1 auto_generated(
	.ram_block3a32(ram_block3a32),
	.ram_block3a0(ram_block3a0),
	.ram_block3a33(ram_block3a33),
	.ram_block3a1(ram_block3a1),
	.ram_block3a34(ram_block3a34),
	.ram_block3a2(ram_block3a2),
	.ram_block3a35(ram_block3a35),
	.ram_block3a3(ram_block3a3),
	.ram_block3a36(ram_block3a36),
	.ram_block3a4(ram_block3a4),
	.ram_block3a37(ram_block3a37),
	.ram_block3a5(ram_block3a5),
	.ram_block3a38(ram_block3a38),
	.ram_block3a6(ram_block3a6),
	.ram_block3a39(ram_block3a39),
	.ram_block3a7(ram_block3a7),
	.ram_block3a40(ram_block3a40),
	.ram_block3a8(ram_block3a8),
	.ram_block3a41(ram_block3a41),
	.ram_block3a9(ram_block3a9),
	.ram_block3a42(ram_block3a42),
	.ram_block3a10(ram_block3a10),
	.ram_block3a43(ram_block3a43),
	.ram_block3a11(ram_block3a11),
	.ram_block3a44(ram_block3a44),
	.ram_block3a12(ram_block3a12),
	.ram_block3a45(ram_block3a45),
	.ram_block3a13(ram_block3a13),
	.ram_block3a46(ram_block3a46),
	.ram_block3a14(ram_block3a14),
	.ram_block3a47(ram_block3a47),
	.ram_block3a15(ram_block3a15),
	.ram_block3a48(ram_block3a48),
	.ram_block3a16(ram_block3a16),
	.ram_block3a49(ram_block3a49),
	.ram_block3a17(ram_block3a17),
	.ram_block3a50(ram_block3a50),
	.ram_block3a18(ram_block3a18),
	.ram_block3a51(ram_block3a51),
	.ram_block3a19(ram_block3a19),
	.ram_block3a52(ram_block3a52),
	.ram_block3a20(ram_block3a20),
	.ram_block3a53(ram_block3a53),
	.ram_block3a21(ram_block3a21),
	.ram_block3a54(ram_block3a54),
	.ram_block3a22(ram_block3a22),
	.ram_block3a55(ram_block3a55),
	.ram_block3a23(ram_block3a23),
	.ram_block3a56(ram_block3a56),
	.ram_block3a24(ram_block3a24),
	.ram_block3a57(ram_block3a57),
	.ram_block3a25(ram_block3a25),
	.ram_block3a58(ram_block3a58),
	.ram_block3a26(ram_block3a26),
	.ram_block3a59(ram_block3a59),
	.ram_block3a27(ram_block3a27),
	.ram_block3a60(ram_block3a60),
	.ram_block3a28(ram_block3a28),
	.ram_block3a61(ram_block3a61),
	.ram_block3a29(ram_block3a29),
	.ram_block3a62(ram_block3a62),
	.ram_block3a30(ram_block3a30),
	.ram_block3a63(ram_block3a63),
	.ram_block3a31(ram_block3a31),
	.is_in_use_reg(is_in_use_reg),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.ramaddr1(ramaddr1),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.irf_reg_0_1(irf_reg_0_1),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_3_1(irf_reg_3_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr_reg(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.altera_internal_jtag1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_99f1 (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	data_a,
	ramaddr1,
	altera_internal_jtag,
	state_4,
	irf_reg_0_1,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_3_1,
	irf_reg_4_1,
	node_ena_1,
	clr_reg,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	altera_internal_jtag1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a32;
output 	ram_block3a0;
output 	ram_block3a33;
output 	ram_block3a1;
output 	ram_block3a34;
output 	ram_block3a2;
output 	ram_block3a35;
output 	ram_block3a3;
output 	ram_block3a36;
output 	ram_block3a4;
output 	ram_block3a37;
output 	ram_block3a5;
output 	ram_block3a38;
output 	ram_block3a6;
output 	ram_block3a39;
output 	ram_block3a7;
output 	ram_block3a40;
output 	ram_block3a8;
output 	ram_block3a41;
output 	ram_block3a9;
output 	ram_block3a42;
output 	ram_block3a10;
output 	ram_block3a43;
output 	ram_block3a11;
output 	ram_block3a44;
output 	ram_block3a12;
output 	ram_block3a45;
output 	ram_block3a13;
output 	ram_block3a46;
output 	ram_block3a14;
output 	ram_block3a47;
output 	ram_block3a15;
output 	ram_block3a48;
output 	ram_block3a16;
output 	ram_block3a49;
output 	ram_block3a17;
output 	ram_block3a50;
output 	ram_block3a18;
output 	ram_block3a51;
output 	ram_block3a19;
output 	ram_block3a52;
output 	ram_block3a20;
output 	ram_block3a53;
output 	ram_block3a21;
output 	ram_block3a54;
output 	ram_block3a22;
output 	ram_block3a55;
output 	ram_block3a23;
output 	ram_block3a56;
output 	ram_block3a24;
output 	ram_block3a57;
output 	ram_block3a25;
output 	ram_block3a58;
output 	ram_block3a26;
output 	ram_block3a59;
output 	ram_block3a27;
output 	ram_block3a60;
output 	ram_block3a28;
output 	ram_block3a61;
output 	ram_block3a29;
output 	ram_block3a62;
output 	ram_block3a30;
output 	ram_block3a63;
output 	ram_block3a31;
output 	is_in_use_reg;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
input 	[31:0] data_a;
input 	ramaddr1;
input 	altera_internal_jtag;
input 	state_4;
input 	irf_reg_0_1;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_3_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr_reg;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	altera_internal_jtag1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \altsyncram1|ram_block3a32~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a0~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a33~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a1~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a34~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a2~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a35~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a3~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a36~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a4~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a37~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a5~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a38~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a6~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a39~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a7~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a40~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a8~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a41~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a9~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a42~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a10~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a43~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a11~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a44~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a12~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a45~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a13~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a46~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a14~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a47~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a15~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a48~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a16~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a49~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a17~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a50~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a18~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a51~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a19~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a52~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a20~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a53~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a21~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a54~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a22~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a55~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a23~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a56~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a24~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a57~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a25~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a58~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a26~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a59~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a27~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a60~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a28~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a61~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a29~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a62~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a30~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a63~PORTBDATAOUT0 ;
wire \altsyncram1|ram_block3a31~PORTBDATAOUT0 ;
wire \mgl_prim2|sdr~0_combout ;
wire [0:0] \altsyncram1|address_reg_b ;
wire [31:0] \mgl_prim2|ram_rom_data_reg ;
wire [13:0] \mgl_prim2|ram_rom_addr_reg ;


sld_mod_ram_rom mgl_prim2(
	.ram_block3a32(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a0(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a33(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a1(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a34(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a2(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a35(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a3(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a36(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a4(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a37(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a5(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a38(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a6(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a39(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a7(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a40(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a8(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a41(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a9(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a42(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a10(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a43(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a11(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a44(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a12(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a45(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a13(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a46(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a14(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a47(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a15(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a48(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a16(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a49(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a17(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a50(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a18(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a51(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a19(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a52(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a20(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a53(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a21(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a54(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a22(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a55(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a23(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a56(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a24(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a57(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a25(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a58(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a26(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a59(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a27(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a60(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a28(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a61(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a29(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a62(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a30(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a63(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a31(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.is_in_use_reg1(is_in_use_reg),
	.ram_rom_data_reg_0(\mgl_prim2|ram_rom_data_reg [0]),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.ram_rom_addr_reg_0(\mgl_prim2|ram_rom_addr_reg [0]),
	.ram_rom_addr_reg_1(\mgl_prim2|ram_rom_addr_reg [1]),
	.ram_rom_addr_reg_2(\mgl_prim2|ram_rom_addr_reg [2]),
	.ram_rom_addr_reg_3(\mgl_prim2|ram_rom_addr_reg [3]),
	.ram_rom_addr_reg_4(\mgl_prim2|ram_rom_addr_reg [4]),
	.ram_rom_addr_reg_5(\mgl_prim2|ram_rom_addr_reg [5]),
	.ram_rom_addr_reg_6(\mgl_prim2|ram_rom_addr_reg [6]),
	.ram_rom_addr_reg_7(\mgl_prim2|ram_rom_addr_reg [7]),
	.ram_rom_addr_reg_8(\mgl_prim2|ram_rom_addr_reg [8]),
	.ram_rom_addr_reg_9(\mgl_prim2|ram_rom_addr_reg [9]),
	.ram_rom_addr_reg_10(\mgl_prim2|ram_rom_addr_reg [10]),
	.ram_rom_addr_reg_11(\mgl_prim2|ram_rom_addr_reg [11]),
	.ram_rom_addr_reg_12(\mgl_prim2|ram_rom_addr_reg [12]),
	.ram_rom_data_reg_1(\mgl_prim2|ram_rom_data_reg [1]),
	.ram_rom_data_reg_2(\mgl_prim2|ram_rom_data_reg [2]),
	.ram_rom_data_reg_3(\mgl_prim2|ram_rom_data_reg [3]),
	.ram_rom_data_reg_4(\mgl_prim2|ram_rom_data_reg [4]),
	.ram_rom_data_reg_5(\mgl_prim2|ram_rom_data_reg [5]),
	.ram_rom_data_reg_6(\mgl_prim2|ram_rom_data_reg [6]),
	.ram_rom_data_reg_7(\mgl_prim2|ram_rom_data_reg [7]),
	.ram_rom_data_reg_8(\mgl_prim2|ram_rom_data_reg [8]),
	.ram_rom_data_reg_9(\mgl_prim2|ram_rom_data_reg [9]),
	.ram_rom_data_reg_10(\mgl_prim2|ram_rom_data_reg [10]),
	.ram_rom_data_reg_11(\mgl_prim2|ram_rom_data_reg [11]),
	.ram_rom_data_reg_12(\mgl_prim2|ram_rom_data_reg [12]),
	.ram_rom_data_reg_13(\mgl_prim2|ram_rom_data_reg [13]),
	.ram_rom_data_reg_14(\mgl_prim2|ram_rom_data_reg [14]),
	.ram_rom_data_reg_15(\mgl_prim2|ram_rom_data_reg [15]),
	.ram_rom_data_reg_16(\mgl_prim2|ram_rom_data_reg [16]),
	.ram_rom_data_reg_17(\mgl_prim2|ram_rom_data_reg [17]),
	.ram_rom_data_reg_18(\mgl_prim2|ram_rom_data_reg [18]),
	.ram_rom_data_reg_19(\mgl_prim2|ram_rom_data_reg [19]),
	.ram_rom_data_reg_20(\mgl_prim2|ram_rom_data_reg [20]),
	.ram_rom_data_reg_21(\mgl_prim2|ram_rom_data_reg [21]),
	.ram_rom_data_reg_22(\mgl_prim2|ram_rom_data_reg [22]),
	.ram_rom_data_reg_23(\mgl_prim2|ram_rom_data_reg [23]),
	.ram_rom_data_reg_24(\mgl_prim2|ram_rom_data_reg [24]),
	.ram_rom_data_reg_25(\mgl_prim2|ram_rom_data_reg [25]),
	.ram_rom_data_reg_26(\mgl_prim2|ram_rom_data_reg [26]),
	.ram_rom_data_reg_27(\mgl_prim2|ram_rom_data_reg [27]),
	.ram_rom_data_reg_28(\mgl_prim2|ram_rom_data_reg [28]),
	.ram_rom_data_reg_29(\mgl_prim2|ram_rom_data_reg [29]),
	.ram_rom_data_reg_30(\mgl_prim2|ram_rom_data_reg [30]),
	.ram_rom_data_reg_31(\mgl_prim2|ram_rom_data_reg [31]),
	.ir_loaded_address_reg_0(ir_loaded_address_reg_0),
	.ir_loaded_address_reg_1(ir_loaded_address_reg_1),
	.ir_loaded_address_reg_2(ir_loaded_address_reg_2),
	.ir_loaded_address_reg_3(ir_loaded_address_reg_3),
	.tdo(tdo),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.ir_in({gnd,irf_reg_3_1,gnd,gnd,irf_reg_0_1}),
	.irf_reg_1_1(irf_reg_1_1),
	.irf_reg_2_1(irf_reg_2_1),
	.irf_reg_4_1(irf_reg_4_1),
	.node_ena_1(node_ena_1),
	.clr(clr_reg),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_5(state_5),
	.state_8(state_8),
	.raw_tck(altera_internal_jtag1),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

altsyncram_fta2 altsyncram1(
	.ram_block3a321(ram_block3a32),
	.ram_block3a322(\altsyncram1|ram_block3a32~PORTBDATAOUT0 ),
	.ram_block3a01(ram_block3a0),
	.ram_block3a02(\altsyncram1|ram_block3a0~PORTBDATAOUT0 ),
	.ram_block3a331(ram_block3a33),
	.ram_block3a332(\altsyncram1|ram_block3a33~PORTBDATAOUT0 ),
	.ram_block3a110(ram_block3a1),
	.ram_block3a111(\altsyncram1|ram_block3a1~PORTBDATAOUT0 ),
	.ram_block3a341(ram_block3a34),
	.ram_block3a342(\altsyncram1|ram_block3a34~PORTBDATAOUT0 ),
	.ram_block3a210(ram_block3a2),
	.ram_block3a211(\altsyncram1|ram_block3a2~PORTBDATAOUT0 ),
	.ram_block3a351(ram_block3a35),
	.ram_block3a352(\altsyncram1|ram_block3a35~PORTBDATAOUT0 ),
	.ram_block3a310(ram_block3a3),
	.ram_block3a311(\altsyncram1|ram_block3a3~PORTBDATAOUT0 ),
	.ram_block3a361(ram_block3a36),
	.ram_block3a362(\altsyncram1|ram_block3a36~PORTBDATAOUT0 ),
	.ram_block3a410(ram_block3a4),
	.ram_block3a411(\altsyncram1|ram_block3a4~PORTBDATAOUT0 ),
	.ram_block3a371(ram_block3a37),
	.ram_block3a372(\altsyncram1|ram_block3a37~PORTBDATAOUT0 ),
	.ram_block3a510(ram_block3a5),
	.ram_block3a511(\altsyncram1|ram_block3a5~PORTBDATAOUT0 ),
	.ram_block3a381(ram_block3a38),
	.ram_block3a382(\altsyncram1|ram_block3a38~PORTBDATAOUT0 ),
	.ram_block3a64(ram_block3a6),
	.ram_block3a65(\altsyncram1|ram_block3a6~PORTBDATAOUT0 ),
	.ram_block3a391(ram_block3a39),
	.ram_block3a392(\altsyncram1|ram_block3a39~PORTBDATAOUT0 ),
	.ram_block3a71(ram_block3a7),
	.ram_block3a72(\altsyncram1|ram_block3a7~PORTBDATAOUT0 ),
	.ram_block3a401(ram_block3a40),
	.ram_block3a402(\altsyncram1|ram_block3a40~PORTBDATAOUT0 ),
	.ram_block3a81(ram_block3a8),
	.ram_block3a82(\altsyncram1|ram_block3a8~PORTBDATAOUT0 ),
	.ram_block3a412(ram_block3a41),
	.ram_block3a413(\altsyncram1|ram_block3a41~PORTBDATAOUT0 ),
	.ram_block3a91(ram_block3a9),
	.ram_block3a92(\altsyncram1|ram_block3a9~PORTBDATAOUT0 ),
	.ram_block3a421(ram_block3a42),
	.ram_block3a422(\altsyncram1|ram_block3a42~PORTBDATAOUT0 ),
	.ram_block3a101(ram_block3a10),
	.ram_block3a102(\altsyncram1|ram_block3a10~PORTBDATAOUT0 ),
	.ram_block3a431(ram_block3a43),
	.ram_block3a432(\altsyncram1|ram_block3a43~PORTBDATAOUT0 ),
	.ram_block3a112(ram_block3a11),
	.ram_block3a113(\altsyncram1|ram_block3a11~PORTBDATAOUT0 ),
	.ram_block3a441(ram_block3a44),
	.ram_block3a442(\altsyncram1|ram_block3a44~PORTBDATAOUT0 ),
	.ram_block3a121(ram_block3a12),
	.ram_block3a122(\altsyncram1|ram_block3a12~PORTBDATAOUT0 ),
	.ram_block3a451(ram_block3a45),
	.ram_block3a452(\altsyncram1|ram_block3a45~PORTBDATAOUT0 ),
	.ram_block3a131(ram_block3a13),
	.ram_block3a132(\altsyncram1|ram_block3a13~PORTBDATAOUT0 ),
	.ram_block3a461(ram_block3a46),
	.ram_block3a462(\altsyncram1|ram_block3a46~PORTBDATAOUT0 ),
	.ram_block3a141(ram_block3a14),
	.ram_block3a142(\altsyncram1|ram_block3a14~PORTBDATAOUT0 ),
	.ram_block3a471(ram_block3a47),
	.ram_block3a472(\altsyncram1|ram_block3a47~PORTBDATAOUT0 ),
	.ram_block3a151(ram_block3a15),
	.ram_block3a152(\altsyncram1|ram_block3a15~PORTBDATAOUT0 ),
	.ram_block3a481(ram_block3a48),
	.ram_block3a482(\altsyncram1|ram_block3a48~PORTBDATAOUT0 ),
	.ram_block3a161(ram_block3a16),
	.ram_block3a162(\altsyncram1|ram_block3a16~PORTBDATAOUT0 ),
	.ram_block3a491(ram_block3a49),
	.ram_block3a492(\altsyncram1|ram_block3a49~PORTBDATAOUT0 ),
	.ram_block3a171(ram_block3a17),
	.ram_block3a172(\altsyncram1|ram_block3a17~PORTBDATAOUT0 ),
	.ram_block3a501(ram_block3a50),
	.ram_block3a502(\altsyncram1|ram_block3a50~PORTBDATAOUT0 ),
	.ram_block3a181(ram_block3a18),
	.ram_block3a182(\altsyncram1|ram_block3a18~PORTBDATAOUT0 ),
	.ram_block3a512(ram_block3a51),
	.ram_block3a513(\altsyncram1|ram_block3a51~PORTBDATAOUT0 ),
	.ram_block3a191(ram_block3a19),
	.ram_block3a192(\altsyncram1|ram_block3a19~PORTBDATAOUT0 ),
	.ram_block3a521(ram_block3a52),
	.ram_block3a522(\altsyncram1|ram_block3a52~PORTBDATAOUT0 ),
	.ram_block3a201(ram_block3a20),
	.ram_block3a202(\altsyncram1|ram_block3a20~PORTBDATAOUT0 ),
	.ram_block3a531(ram_block3a53),
	.ram_block3a532(\altsyncram1|ram_block3a53~PORTBDATAOUT0 ),
	.ram_block3a212(ram_block3a21),
	.ram_block3a213(\altsyncram1|ram_block3a21~PORTBDATAOUT0 ),
	.ram_block3a541(ram_block3a54),
	.ram_block3a542(\altsyncram1|ram_block3a54~PORTBDATAOUT0 ),
	.ram_block3a221(ram_block3a22),
	.ram_block3a222(\altsyncram1|ram_block3a22~PORTBDATAOUT0 ),
	.ram_block3a551(ram_block3a55),
	.ram_block3a552(\altsyncram1|ram_block3a55~PORTBDATAOUT0 ),
	.ram_block3a231(ram_block3a23),
	.ram_block3a232(\altsyncram1|ram_block3a23~PORTBDATAOUT0 ),
	.ram_block3a561(ram_block3a56),
	.ram_block3a562(\altsyncram1|ram_block3a56~PORTBDATAOUT0 ),
	.ram_block3a241(ram_block3a24),
	.ram_block3a242(\altsyncram1|ram_block3a24~PORTBDATAOUT0 ),
	.ram_block3a571(ram_block3a57),
	.ram_block3a572(\altsyncram1|ram_block3a57~PORTBDATAOUT0 ),
	.ram_block3a251(ram_block3a25),
	.ram_block3a252(\altsyncram1|ram_block3a25~PORTBDATAOUT0 ),
	.ram_block3a581(ram_block3a58),
	.ram_block3a582(\altsyncram1|ram_block3a58~PORTBDATAOUT0 ),
	.ram_block3a261(ram_block3a26),
	.ram_block3a262(\altsyncram1|ram_block3a26~PORTBDATAOUT0 ),
	.ram_block3a591(ram_block3a59),
	.ram_block3a592(\altsyncram1|ram_block3a59~PORTBDATAOUT0 ),
	.ram_block3a271(ram_block3a27),
	.ram_block3a272(\altsyncram1|ram_block3a27~PORTBDATAOUT0 ),
	.ram_block3a601(ram_block3a60),
	.ram_block3a602(\altsyncram1|ram_block3a60~PORTBDATAOUT0 ),
	.ram_block3a281(ram_block3a28),
	.ram_block3a282(\altsyncram1|ram_block3a28~PORTBDATAOUT0 ),
	.ram_block3a611(ram_block3a61),
	.ram_block3a612(\altsyncram1|ram_block3a61~PORTBDATAOUT0 ),
	.ram_block3a291(ram_block3a29),
	.ram_block3a292(\altsyncram1|ram_block3a29~PORTBDATAOUT0 ),
	.ram_block3a621(ram_block3a62),
	.ram_block3a622(\altsyncram1|ram_block3a62~PORTBDATAOUT0 ),
	.ram_block3a301(ram_block3a30),
	.ram_block3a302(\altsyncram1|ram_block3a30~PORTBDATAOUT0 ),
	.ram_block3a631(ram_block3a63),
	.ram_block3a632(\altsyncram1|ram_block3a63~PORTBDATAOUT0 ),
	.ram_block3a312(ram_block3a31),
	.ram_block3a313(\altsyncram1|ram_block3a31~PORTBDATAOUT0 ),
	.data_b({\mgl_prim2|ram_rom_data_reg [31],\mgl_prim2|ram_rom_data_reg [30],\mgl_prim2|ram_rom_data_reg [29],\mgl_prim2|ram_rom_data_reg [28],\mgl_prim2|ram_rom_data_reg [27],\mgl_prim2|ram_rom_data_reg [26],\mgl_prim2|ram_rom_data_reg [25],\mgl_prim2|ram_rom_data_reg [24],\mgl_prim2|ram_rom_data_reg [23],
\mgl_prim2|ram_rom_data_reg [22],\mgl_prim2|ram_rom_data_reg [21],\mgl_prim2|ram_rom_data_reg [20],\mgl_prim2|ram_rom_data_reg [19],\mgl_prim2|ram_rom_data_reg [18],\mgl_prim2|ram_rom_data_reg [17],\mgl_prim2|ram_rom_data_reg [16],\mgl_prim2|ram_rom_data_reg [15],\mgl_prim2|ram_rom_data_reg [14],
\mgl_prim2|ram_rom_data_reg [13],\mgl_prim2|ram_rom_data_reg [12],\mgl_prim2|ram_rom_data_reg [11],\mgl_prim2|ram_rom_data_reg [10],\mgl_prim2|ram_rom_data_reg [9],\mgl_prim2|ram_rom_data_reg [8],\mgl_prim2|ram_rom_data_reg [7],\mgl_prim2|ram_rom_data_reg [6],\mgl_prim2|ram_rom_data_reg [5],
\mgl_prim2|ram_rom_data_reg [4],\mgl_prim2|ram_rom_data_reg [3],\mgl_prim2|ram_rom_data_reg [2],\mgl_prim2|ram_rom_data_reg [1],\mgl_prim2|ram_rom_data_reg [0]}),
	.ram_rom_addr_reg_13(\mgl_prim2|ram_rom_addr_reg [13]),
	.address_b({gnd,\mgl_prim2|ram_rom_addr_reg [12],\mgl_prim2|ram_rom_addr_reg [11],\mgl_prim2|ram_rom_addr_reg [10],\mgl_prim2|ram_rom_addr_reg [9],\mgl_prim2|ram_rom_addr_reg [8],\mgl_prim2|ram_rom_addr_reg [7],\mgl_prim2|ram_rom_addr_reg [6],\mgl_prim2|ram_rom_addr_reg [5],\mgl_prim2|ram_rom_addr_reg [4],
\mgl_prim2|ram_rom_addr_reg [3],\mgl_prim2|ram_rom_addr_reg [2],\mgl_prim2|ram_rom_addr_reg [1],\mgl_prim2|ram_rom_addr_reg [0]}),
	.address_reg_a_0(address_reg_a_0),
	.address_a({gnd,address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.sdr(\mgl_prim2|sdr~0_combout ),
	.data_a({data_a[31],data_a[30],data_a[29],data_a[28],data_a[27],data_a[26],data_a[25],data_a[24],data_a[23],data_a[22],data_a[21],data_a[20],data_a[19],data_a[18],data_a[17],data_a[16],data_a[15],data_a[14],data_a[13],data_a[12],data_a[11],data_a[10],data_a[9],data_a[8],data_a[7],data_a[6],data_a[5],data_a[4],data_a[3],data_a[2],data_a[1],data_a[0]}),
	.address_reg_b_0(\altsyncram1|address_reg_b [0]),
	.ramaddr1(ramaddr1),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.clock1(altera_internal_jtag1),
	.clock0(clock0),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

endmodule

module altsyncram_fta2 (
	ram_block3a321,
	ram_block3a322,
	ram_block3a01,
	ram_block3a02,
	ram_block3a331,
	ram_block3a332,
	ram_block3a110,
	ram_block3a111,
	ram_block3a341,
	ram_block3a342,
	ram_block3a210,
	ram_block3a211,
	ram_block3a351,
	ram_block3a352,
	ram_block3a310,
	ram_block3a311,
	ram_block3a361,
	ram_block3a362,
	ram_block3a410,
	ram_block3a411,
	ram_block3a371,
	ram_block3a372,
	ram_block3a510,
	ram_block3a511,
	ram_block3a381,
	ram_block3a382,
	ram_block3a64,
	ram_block3a65,
	ram_block3a391,
	ram_block3a392,
	ram_block3a71,
	ram_block3a72,
	ram_block3a401,
	ram_block3a402,
	ram_block3a81,
	ram_block3a82,
	ram_block3a412,
	ram_block3a413,
	ram_block3a91,
	ram_block3a92,
	ram_block3a421,
	ram_block3a422,
	ram_block3a101,
	ram_block3a102,
	ram_block3a431,
	ram_block3a432,
	ram_block3a112,
	ram_block3a113,
	ram_block3a441,
	ram_block3a442,
	ram_block3a121,
	ram_block3a122,
	ram_block3a451,
	ram_block3a452,
	ram_block3a131,
	ram_block3a132,
	ram_block3a461,
	ram_block3a462,
	ram_block3a141,
	ram_block3a142,
	ram_block3a471,
	ram_block3a472,
	ram_block3a151,
	ram_block3a152,
	ram_block3a481,
	ram_block3a482,
	ram_block3a161,
	ram_block3a162,
	ram_block3a491,
	ram_block3a492,
	ram_block3a171,
	ram_block3a172,
	ram_block3a501,
	ram_block3a502,
	ram_block3a181,
	ram_block3a182,
	ram_block3a512,
	ram_block3a513,
	ram_block3a191,
	ram_block3a192,
	ram_block3a521,
	ram_block3a522,
	ram_block3a201,
	ram_block3a202,
	ram_block3a531,
	ram_block3a532,
	ram_block3a212,
	ram_block3a213,
	ram_block3a541,
	ram_block3a542,
	ram_block3a221,
	ram_block3a222,
	ram_block3a551,
	ram_block3a552,
	ram_block3a231,
	ram_block3a232,
	ram_block3a561,
	ram_block3a562,
	ram_block3a241,
	ram_block3a242,
	ram_block3a571,
	ram_block3a572,
	ram_block3a251,
	ram_block3a252,
	ram_block3a581,
	ram_block3a582,
	ram_block3a261,
	ram_block3a262,
	ram_block3a591,
	ram_block3a592,
	ram_block3a271,
	ram_block3a272,
	ram_block3a601,
	ram_block3a602,
	ram_block3a281,
	ram_block3a282,
	ram_block3a611,
	ram_block3a612,
	ram_block3a291,
	ram_block3a292,
	ram_block3a621,
	ram_block3a622,
	ram_block3a301,
	ram_block3a302,
	ram_block3a631,
	ram_block3a632,
	ram_block3a312,
	ram_block3a313,
	data_b,
	ram_rom_addr_reg_13,
	address_b,
	address_reg_a_0,
	address_a,
	ramaddr,
	ramWEN,
	always1,
	sdr,
	data_a,
	address_reg_b_0,
	ramaddr1,
	irf_reg_2_1,
	state_5,
	clock1,
	clock0,
	devpor,
	devclrn,
	devoe);
output 	ram_block3a321;
output 	ram_block3a322;
output 	ram_block3a01;
output 	ram_block3a02;
output 	ram_block3a331;
output 	ram_block3a332;
output 	ram_block3a110;
output 	ram_block3a111;
output 	ram_block3a341;
output 	ram_block3a342;
output 	ram_block3a210;
output 	ram_block3a211;
output 	ram_block3a351;
output 	ram_block3a352;
output 	ram_block3a310;
output 	ram_block3a311;
output 	ram_block3a361;
output 	ram_block3a362;
output 	ram_block3a410;
output 	ram_block3a411;
output 	ram_block3a371;
output 	ram_block3a372;
output 	ram_block3a510;
output 	ram_block3a511;
output 	ram_block3a381;
output 	ram_block3a382;
output 	ram_block3a64;
output 	ram_block3a65;
output 	ram_block3a391;
output 	ram_block3a392;
output 	ram_block3a71;
output 	ram_block3a72;
output 	ram_block3a401;
output 	ram_block3a402;
output 	ram_block3a81;
output 	ram_block3a82;
output 	ram_block3a412;
output 	ram_block3a413;
output 	ram_block3a91;
output 	ram_block3a92;
output 	ram_block3a421;
output 	ram_block3a422;
output 	ram_block3a101;
output 	ram_block3a102;
output 	ram_block3a431;
output 	ram_block3a432;
output 	ram_block3a112;
output 	ram_block3a113;
output 	ram_block3a441;
output 	ram_block3a442;
output 	ram_block3a121;
output 	ram_block3a122;
output 	ram_block3a451;
output 	ram_block3a452;
output 	ram_block3a131;
output 	ram_block3a132;
output 	ram_block3a461;
output 	ram_block3a462;
output 	ram_block3a141;
output 	ram_block3a142;
output 	ram_block3a471;
output 	ram_block3a472;
output 	ram_block3a151;
output 	ram_block3a152;
output 	ram_block3a481;
output 	ram_block3a482;
output 	ram_block3a161;
output 	ram_block3a162;
output 	ram_block3a491;
output 	ram_block3a492;
output 	ram_block3a171;
output 	ram_block3a172;
output 	ram_block3a501;
output 	ram_block3a502;
output 	ram_block3a181;
output 	ram_block3a182;
output 	ram_block3a512;
output 	ram_block3a513;
output 	ram_block3a191;
output 	ram_block3a192;
output 	ram_block3a521;
output 	ram_block3a522;
output 	ram_block3a201;
output 	ram_block3a202;
output 	ram_block3a531;
output 	ram_block3a532;
output 	ram_block3a212;
output 	ram_block3a213;
output 	ram_block3a541;
output 	ram_block3a542;
output 	ram_block3a221;
output 	ram_block3a222;
output 	ram_block3a551;
output 	ram_block3a552;
output 	ram_block3a231;
output 	ram_block3a232;
output 	ram_block3a561;
output 	ram_block3a562;
output 	ram_block3a241;
output 	ram_block3a242;
output 	ram_block3a571;
output 	ram_block3a572;
output 	ram_block3a251;
output 	ram_block3a252;
output 	ram_block3a581;
output 	ram_block3a582;
output 	ram_block3a261;
output 	ram_block3a262;
output 	ram_block3a591;
output 	ram_block3a592;
output 	ram_block3a271;
output 	ram_block3a272;
output 	ram_block3a601;
output 	ram_block3a602;
output 	ram_block3a281;
output 	ram_block3a282;
output 	ram_block3a611;
output 	ram_block3a612;
output 	ram_block3a291;
output 	ram_block3a292;
output 	ram_block3a621;
output 	ram_block3a622;
output 	ram_block3a301;
output 	ram_block3a302;
output 	ram_block3a631;
output 	ram_block3a632;
output 	ram_block3a312;
output 	ram_block3a313;
input 	[31:0] data_b;
input 	ram_rom_addr_reg_13;
input 	[13:0] address_b;
output 	address_reg_a_0;
input 	[13:0] address_a;
input 	ramaddr;
input 	ramWEN;
input 	always1;
input 	sdr;
input 	[31:0] data_a;
output 	address_reg_b_0;
input 	ramaddr1;
input 	irf_reg_2_1;
input 	state_5;
input 	clock1;
input 	clock0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \decode4|eq_node[1]~0_combout ;
wire \decode5|eq_node[1]~0_combout ;
wire \decode4|eq_node[0]~1_combout ;
wire \decode5|eq_node[0]~1_combout ;
wire \address_reg_b[0]~feeder_combout ;

wire [0:0] ram_block3a32_PORTADATAOUT_bus;
wire [0:0] ram_block3a32_PORTBDATAOUT_bus;
wire [0:0] ram_block3a0_PORTADATAOUT_bus;
wire [0:0] ram_block3a0_PORTBDATAOUT_bus;
wire [0:0] ram_block3a33_PORTADATAOUT_bus;
wire [0:0] ram_block3a33_PORTBDATAOUT_bus;
wire [0:0] ram_block3a1_PORTADATAOUT_bus;
wire [0:0] ram_block3a1_PORTBDATAOUT_bus;
wire [0:0] ram_block3a34_PORTADATAOUT_bus;
wire [0:0] ram_block3a34_PORTBDATAOUT_bus;
wire [0:0] ram_block3a2_PORTADATAOUT_bus;
wire [0:0] ram_block3a2_PORTBDATAOUT_bus;
wire [0:0] ram_block3a35_PORTADATAOUT_bus;
wire [0:0] ram_block3a35_PORTBDATAOUT_bus;
wire [0:0] ram_block3a3_PORTADATAOUT_bus;
wire [0:0] ram_block3a3_PORTBDATAOUT_bus;
wire [0:0] ram_block3a36_PORTADATAOUT_bus;
wire [0:0] ram_block3a36_PORTBDATAOUT_bus;
wire [0:0] ram_block3a4_PORTADATAOUT_bus;
wire [0:0] ram_block3a4_PORTBDATAOUT_bus;
wire [0:0] ram_block3a37_PORTADATAOUT_bus;
wire [0:0] ram_block3a37_PORTBDATAOUT_bus;
wire [0:0] ram_block3a5_PORTADATAOUT_bus;
wire [0:0] ram_block3a5_PORTBDATAOUT_bus;
wire [0:0] ram_block3a38_PORTADATAOUT_bus;
wire [0:0] ram_block3a38_PORTBDATAOUT_bus;
wire [0:0] ram_block3a6_PORTADATAOUT_bus;
wire [0:0] ram_block3a6_PORTBDATAOUT_bus;
wire [0:0] ram_block3a39_PORTADATAOUT_bus;
wire [0:0] ram_block3a39_PORTBDATAOUT_bus;
wire [0:0] ram_block3a7_PORTADATAOUT_bus;
wire [0:0] ram_block3a7_PORTBDATAOUT_bus;
wire [0:0] ram_block3a40_PORTADATAOUT_bus;
wire [0:0] ram_block3a40_PORTBDATAOUT_bus;
wire [0:0] ram_block3a8_PORTADATAOUT_bus;
wire [0:0] ram_block3a8_PORTBDATAOUT_bus;
wire [0:0] ram_block3a41_PORTADATAOUT_bus;
wire [0:0] ram_block3a41_PORTBDATAOUT_bus;
wire [0:0] ram_block3a9_PORTADATAOUT_bus;
wire [0:0] ram_block3a9_PORTBDATAOUT_bus;
wire [0:0] ram_block3a42_PORTADATAOUT_bus;
wire [0:0] ram_block3a42_PORTBDATAOUT_bus;
wire [0:0] ram_block3a10_PORTADATAOUT_bus;
wire [0:0] ram_block3a10_PORTBDATAOUT_bus;
wire [0:0] ram_block3a43_PORTADATAOUT_bus;
wire [0:0] ram_block3a43_PORTBDATAOUT_bus;
wire [0:0] ram_block3a11_PORTADATAOUT_bus;
wire [0:0] ram_block3a11_PORTBDATAOUT_bus;
wire [0:0] ram_block3a44_PORTADATAOUT_bus;
wire [0:0] ram_block3a44_PORTBDATAOUT_bus;
wire [0:0] ram_block3a12_PORTADATAOUT_bus;
wire [0:0] ram_block3a12_PORTBDATAOUT_bus;
wire [0:0] ram_block3a45_PORTADATAOUT_bus;
wire [0:0] ram_block3a45_PORTBDATAOUT_bus;
wire [0:0] ram_block3a13_PORTADATAOUT_bus;
wire [0:0] ram_block3a13_PORTBDATAOUT_bus;
wire [0:0] ram_block3a46_PORTADATAOUT_bus;
wire [0:0] ram_block3a46_PORTBDATAOUT_bus;
wire [0:0] ram_block3a14_PORTADATAOUT_bus;
wire [0:0] ram_block3a14_PORTBDATAOUT_bus;
wire [0:0] ram_block3a47_PORTADATAOUT_bus;
wire [0:0] ram_block3a47_PORTBDATAOUT_bus;
wire [0:0] ram_block3a15_PORTADATAOUT_bus;
wire [0:0] ram_block3a15_PORTBDATAOUT_bus;
wire [0:0] ram_block3a48_PORTADATAOUT_bus;
wire [0:0] ram_block3a48_PORTBDATAOUT_bus;
wire [0:0] ram_block3a16_PORTADATAOUT_bus;
wire [0:0] ram_block3a16_PORTBDATAOUT_bus;
wire [0:0] ram_block3a49_PORTADATAOUT_bus;
wire [0:0] ram_block3a49_PORTBDATAOUT_bus;
wire [0:0] ram_block3a17_PORTADATAOUT_bus;
wire [0:0] ram_block3a17_PORTBDATAOUT_bus;
wire [0:0] ram_block3a50_PORTADATAOUT_bus;
wire [0:0] ram_block3a50_PORTBDATAOUT_bus;
wire [0:0] ram_block3a18_PORTADATAOUT_bus;
wire [0:0] ram_block3a18_PORTBDATAOUT_bus;
wire [0:0] ram_block3a51_PORTADATAOUT_bus;
wire [0:0] ram_block3a51_PORTBDATAOUT_bus;
wire [0:0] ram_block3a19_PORTADATAOUT_bus;
wire [0:0] ram_block3a19_PORTBDATAOUT_bus;
wire [0:0] ram_block3a52_PORTADATAOUT_bus;
wire [0:0] ram_block3a52_PORTBDATAOUT_bus;
wire [0:0] ram_block3a20_PORTADATAOUT_bus;
wire [0:0] ram_block3a20_PORTBDATAOUT_bus;
wire [0:0] ram_block3a53_PORTADATAOUT_bus;
wire [0:0] ram_block3a53_PORTBDATAOUT_bus;
wire [0:0] ram_block3a21_PORTADATAOUT_bus;
wire [0:0] ram_block3a21_PORTBDATAOUT_bus;
wire [0:0] ram_block3a54_PORTADATAOUT_bus;
wire [0:0] ram_block3a54_PORTBDATAOUT_bus;
wire [0:0] ram_block3a22_PORTADATAOUT_bus;
wire [0:0] ram_block3a22_PORTBDATAOUT_bus;
wire [0:0] ram_block3a55_PORTADATAOUT_bus;
wire [0:0] ram_block3a55_PORTBDATAOUT_bus;
wire [0:0] ram_block3a23_PORTADATAOUT_bus;
wire [0:0] ram_block3a23_PORTBDATAOUT_bus;
wire [0:0] ram_block3a56_PORTADATAOUT_bus;
wire [0:0] ram_block3a56_PORTBDATAOUT_bus;
wire [0:0] ram_block3a24_PORTADATAOUT_bus;
wire [0:0] ram_block3a24_PORTBDATAOUT_bus;
wire [0:0] ram_block3a57_PORTADATAOUT_bus;
wire [0:0] ram_block3a57_PORTBDATAOUT_bus;
wire [0:0] ram_block3a25_PORTADATAOUT_bus;
wire [0:0] ram_block3a25_PORTBDATAOUT_bus;
wire [0:0] ram_block3a58_PORTADATAOUT_bus;
wire [0:0] ram_block3a58_PORTBDATAOUT_bus;
wire [0:0] ram_block3a26_PORTADATAOUT_bus;
wire [0:0] ram_block3a26_PORTBDATAOUT_bus;
wire [0:0] ram_block3a59_PORTADATAOUT_bus;
wire [0:0] ram_block3a59_PORTBDATAOUT_bus;
wire [0:0] ram_block3a27_PORTADATAOUT_bus;
wire [0:0] ram_block3a27_PORTBDATAOUT_bus;
wire [0:0] ram_block3a60_PORTADATAOUT_bus;
wire [0:0] ram_block3a60_PORTBDATAOUT_bus;
wire [0:0] ram_block3a28_PORTADATAOUT_bus;
wire [0:0] ram_block3a28_PORTBDATAOUT_bus;
wire [0:0] ram_block3a61_PORTADATAOUT_bus;
wire [0:0] ram_block3a61_PORTBDATAOUT_bus;
wire [0:0] ram_block3a29_PORTADATAOUT_bus;
wire [0:0] ram_block3a29_PORTBDATAOUT_bus;
wire [0:0] ram_block3a62_PORTADATAOUT_bus;
wire [0:0] ram_block3a62_PORTBDATAOUT_bus;
wire [0:0] ram_block3a30_PORTADATAOUT_bus;
wire [0:0] ram_block3a30_PORTBDATAOUT_bus;
wire [0:0] ram_block3a63_PORTADATAOUT_bus;
wire [0:0] ram_block3a63_PORTBDATAOUT_bus;
wire [0:0] ram_block3a31_PORTADATAOUT_bus;
wire [0:0] ram_block3a31_PORTBDATAOUT_bus;

assign ram_block3a321 = ram_block3a32_PORTADATAOUT_bus[0];

assign ram_block3a322 = ram_block3a32_PORTBDATAOUT_bus[0];

assign ram_block3a01 = ram_block3a0_PORTADATAOUT_bus[0];

assign ram_block3a02 = ram_block3a0_PORTBDATAOUT_bus[0];

assign ram_block3a331 = ram_block3a33_PORTADATAOUT_bus[0];

assign ram_block3a332 = ram_block3a33_PORTBDATAOUT_bus[0];

assign ram_block3a110 = ram_block3a1_PORTADATAOUT_bus[0];

assign ram_block3a111 = ram_block3a1_PORTBDATAOUT_bus[0];

assign ram_block3a341 = ram_block3a34_PORTADATAOUT_bus[0];

assign ram_block3a342 = ram_block3a34_PORTBDATAOUT_bus[0];

assign ram_block3a210 = ram_block3a2_PORTADATAOUT_bus[0];

assign ram_block3a211 = ram_block3a2_PORTBDATAOUT_bus[0];

assign ram_block3a351 = ram_block3a35_PORTADATAOUT_bus[0];

assign ram_block3a352 = ram_block3a35_PORTBDATAOUT_bus[0];

assign ram_block3a310 = ram_block3a3_PORTADATAOUT_bus[0];

assign ram_block3a311 = ram_block3a3_PORTBDATAOUT_bus[0];

assign ram_block3a361 = ram_block3a36_PORTADATAOUT_bus[0];

assign ram_block3a362 = ram_block3a36_PORTBDATAOUT_bus[0];

assign ram_block3a410 = ram_block3a4_PORTADATAOUT_bus[0];

assign ram_block3a411 = ram_block3a4_PORTBDATAOUT_bus[0];

assign ram_block3a371 = ram_block3a37_PORTADATAOUT_bus[0];

assign ram_block3a372 = ram_block3a37_PORTBDATAOUT_bus[0];

assign ram_block3a510 = ram_block3a5_PORTADATAOUT_bus[0];

assign ram_block3a511 = ram_block3a5_PORTBDATAOUT_bus[0];

assign ram_block3a381 = ram_block3a38_PORTADATAOUT_bus[0];

assign ram_block3a382 = ram_block3a38_PORTBDATAOUT_bus[0];

assign ram_block3a64 = ram_block3a6_PORTADATAOUT_bus[0];

assign ram_block3a65 = ram_block3a6_PORTBDATAOUT_bus[0];

assign ram_block3a391 = ram_block3a39_PORTADATAOUT_bus[0];

assign ram_block3a392 = ram_block3a39_PORTBDATAOUT_bus[0];

assign ram_block3a71 = ram_block3a7_PORTADATAOUT_bus[0];

assign ram_block3a72 = ram_block3a7_PORTBDATAOUT_bus[0];

assign ram_block3a401 = ram_block3a40_PORTADATAOUT_bus[0];

assign ram_block3a402 = ram_block3a40_PORTBDATAOUT_bus[0];

assign ram_block3a81 = ram_block3a8_PORTADATAOUT_bus[0];

assign ram_block3a82 = ram_block3a8_PORTBDATAOUT_bus[0];

assign ram_block3a412 = ram_block3a41_PORTADATAOUT_bus[0];

assign ram_block3a413 = ram_block3a41_PORTBDATAOUT_bus[0];

assign ram_block3a91 = ram_block3a9_PORTADATAOUT_bus[0];

assign ram_block3a92 = ram_block3a9_PORTBDATAOUT_bus[0];

assign ram_block3a421 = ram_block3a42_PORTADATAOUT_bus[0];

assign ram_block3a422 = ram_block3a42_PORTBDATAOUT_bus[0];

assign ram_block3a101 = ram_block3a10_PORTADATAOUT_bus[0];

assign ram_block3a102 = ram_block3a10_PORTBDATAOUT_bus[0];

assign ram_block3a431 = ram_block3a43_PORTADATAOUT_bus[0];

assign ram_block3a432 = ram_block3a43_PORTBDATAOUT_bus[0];

assign ram_block3a112 = ram_block3a11_PORTADATAOUT_bus[0];

assign ram_block3a113 = ram_block3a11_PORTBDATAOUT_bus[0];

assign ram_block3a441 = ram_block3a44_PORTADATAOUT_bus[0];

assign ram_block3a442 = ram_block3a44_PORTBDATAOUT_bus[0];

assign ram_block3a121 = ram_block3a12_PORTADATAOUT_bus[0];

assign ram_block3a122 = ram_block3a12_PORTBDATAOUT_bus[0];

assign ram_block3a451 = ram_block3a45_PORTADATAOUT_bus[0];

assign ram_block3a452 = ram_block3a45_PORTBDATAOUT_bus[0];

assign ram_block3a131 = ram_block3a13_PORTADATAOUT_bus[0];

assign ram_block3a132 = ram_block3a13_PORTBDATAOUT_bus[0];

assign ram_block3a461 = ram_block3a46_PORTADATAOUT_bus[0];

assign ram_block3a462 = ram_block3a46_PORTBDATAOUT_bus[0];

assign ram_block3a141 = ram_block3a14_PORTADATAOUT_bus[0];

assign ram_block3a142 = ram_block3a14_PORTBDATAOUT_bus[0];

assign ram_block3a471 = ram_block3a47_PORTADATAOUT_bus[0];

assign ram_block3a472 = ram_block3a47_PORTBDATAOUT_bus[0];

assign ram_block3a151 = ram_block3a15_PORTADATAOUT_bus[0];

assign ram_block3a152 = ram_block3a15_PORTBDATAOUT_bus[0];

assign ram_block3a481 = ram_block3a48_PORTADATAOUT_bus[0];

assign ram_block3a482 = ram_block3a48_PORTBDATAOUT_bus[0];

assign ram_block3a161 = ram_block3a16_PORTADATAOUT_bus[0];

assign ram_block3a162 = ram_block3a16_PORTBDATAOUT_bus[0];

assign ram_block3a491 = ram_block3a49_PORTADATAOUT_bus[0];

assign ram_block3a492 = ram_block3a49_PORTBDATAOUT_bus[0];

assign ram_block3a171 = ram_block3a17_PORTADATAOUT_bus[0];

assign ram_block3a172 = ram_block3a17_PORTBDATAOUT_bus[0];

assign ram_block3a501 = ram_block3a50_PORTADATAOUT_bus[0];

assign ram_block3a502 = ram_block3a50_PORTBDATAOUT_bus[0];

assign ram_block3a181 = ram_block3a18_PORTADATAOUT_bus[0];

assign ram_block3a182 = ram_block3a18_PORTBDATAOUT_bus[0];

assign ram_block3a512 = ram_block3a51_PORTADATAOUT_bus[0];

assign ram_block3a513 = ram_block3a51_PORTBDATAOUT_bus[0];

assign ram_block3a191 = ram_block3a19_PORTADATAOUT_bus[0];

assign ram_block3a192 = ram_block3a19_PORTBDATAOUT_bus[0];

assign ram_block3a521 = ram_block3a52_PORTADATAOUT_bus[0];

assign ram_block3a522 = ram_block3a52_PORTBDATAOUT_bus[0];

assign ram_block3a201 = ram_block3a20_PORTADATAOUT_bus[0];

assign ram_block3a202 = ram_block3a20_PORTBDATAOUT_bus[0];

assign ram_block3a531 = ram_block3a53_PORTADATAOUT_bus[0];

assign ram_block3a532 = ram_block3a53_PORTBDATAOUT_bus[0];

assign ram_block3a212 = ram_block3a21_PORTADATAOUT_bus[0];

assign ram_block3a213 = ram_block3a21_PORTBDATAOUT_bus[0];

assign ram_block3a541 = ram_block3a54_PORTADATAOUT_bus[0];

assign ram_block3a542 = ram_block3a54_PORTBDATAOUT_bus[0];

assign ram_block3a221 = ram_block3a22_PORTADATAOUT_bus[0];

assign ram_block3a222 = ram_block3a22_PORTBDATAOUT_bus[0];

assign ram_block3a551 = ram_block3a55_PORTADATAOUT_bus[0];

assign ram_block3a552 = ram_block3a55_PORTBDATAOUT_bus[0];

assign ram_block3a231 = ram_block3a23_PORTADATAOUT_bus[0];

assign ram_block3a232 = ram_block3a23_PORTBDATAOUT_bus[0];

assign ram_block3a561 = ram_block3a56_PORTADATAOUT_bus[0];

assign ram_block3a562 = ram_block3a56_PORTBDATAOUT_bus[0];

assign ram_block3a241 = ram_block3a24_PORTADATAOUT_bus[0];

assign ram_block3a242 = ram_block3a24_PORTBDATAOUT_bus[0];

assign ram_block3a571 = ram_block3a57_PORTADATAOUT_bus[0];

assign ram_block3a572 = ram_block3a57_PORTBDATAOUT_bus[0];

assign ram_block3a251 = ram_block3a25_PORTADATAOUT_bus[0];

assign ram_block3a252 = ram_block3a25_PORTBDATAOUT_bus[0];

assign ram_block3a581 = ram_block3a58_PORTADATAOUT_bus[0];

assign ram_block3a582 = ram_block3a58_PORTBDATAOUT_bus[0];

assign ram_block3a261 = ram_block3a26_PORTADATAOUT_bus[0];

assign ram_block3a262 = ram_block3a26_PORTBDATAOUT_bus[0];

assign ram_block3a591 = ram_block3a59_PORTADATAOUT_bus[0];

assign ram_block3a592 = ram_block3a59_PORTBDATAOUT_bus[0];

assign ram_block3a271 = ram_block3a27_PORTADATAOUT_bus[0];

assign ram_block3a272 = ram_block3a27_PORTBDATAOUT_bus[0];

assign ram_block3a601 = ram_block3a60_PORTADATAOUT_bus[0];

assign ram_block3a602 = ram_block3a60_PORTBDATAOUT_bus[0];

assign ram_block3a281 = ram_block3a28_PORTADATAOUT_bus[0];

assign ram_block3a282 = ram_block3a28_PORTBDATAOUT_bus[0];

assign ram_block3a611 = ram_block3a61_PORTADATAOUT_bus[0];

assign ram_block3a612 = ram_block3a61_PORTBDATAOUT_bus[0];

assign ram_block3a291 = ram_block3a29_PORTADATAOUT_bus[0];

assign ram_block3a292 = ram_block3a29_PORTBDATAOUT_bus[0];

assign ram_block3a621 = ram_block3a62_PORTADATAOUT_bus[0];

assign ram_block3a622 = ram_block3a62_PORTBDATAOUT_bus[0];

assign ram_block3a301 = ram_block3a30_PORTADATAOUT_bus[0];

assign ram_block3a302 = ram_block3a30_PORTBDATAOUT_bus[0];

assign ram_block3a631 = ram_block3a63_PORTADATAOUT_bus[0];

assign ram_block3a632 = ram_block3a63_PORTBDATAOUT_bus[0];

assign ram_block3a312 = ram_block3a31_PORTADATAOUT_bus[0];

assign ram_block3a313 = ram_block3a31_PORTBDATAOUT_bus[0];

decode_jsa_1 decode5(
	.ram_rom_addr_reg_13(ram_rom_addr_reg_13),
	.sdr(sdr),
	.eq_node_1(\decode5|eq_node[1]~0_combout ),
	.eq_node_0(\decode5|eq_node[0]~1_combout ),
	.irf_reg_2_1(irf_reg_2_1),
	.state_5(state_5),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

decode_jsa decode4(
	.ramaddr(ramaddr),
	.ramWEN(ramWEN),
	.always1(always1),
	.eq_node_1(\decode4|eq_node[1]~0_combout ),
	.eq_node_0(\decode4|eq_node[0]~1_combout ),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: M9K_X51_Y29_N0
cycloneive_ram_block ram_block3a32(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a32_PORTADATAOUT_bus),
	.portbdataout(ram_block3a32_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a32.clk0_core_clock_enable = "ena0";
defparam ram_block3a32.clk1_core_clock_enable = "ena1";
defparam ram_block3a32.data_interleave_offset_in_bits = 1;
defparam ram_block3a32.data_interleave_width_in_bits = 1;
defparam ram_block3a32.init_file = "meminit.hex";
defparam ram_block3a32.init_file_layout = "port_a";
defparam ram_block3a32.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a32.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a32.operation_mode = "bidir_dual_port";
defparam ram_block3a32.port_a_address_clear = "none";
defparam ram_block3a32.port_a_address_width = 13;
defparam ram_block3a32.port_a_byte_enable_clock = "none";
defparam ram_block3a32.port_a_data_out_clear = "none";
defparam ram_block3a32.port_a_data_out_clock = "none";
defparam ram_block3a32.port_a_data_width = 1;
defparam ram_block3a32.port_a_first_address = 0;
defparam ram_block3a32.port_a_first_bit_number = 0;
defparam ram_block3a32.port_a_last_address = 8191;
defparam ram_block3a32.port_a_logical_ram_depth = 16384;
defparam ram_block3a32.port_a_logical_ram_width = 32;
defparam ram_block3a32.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_address_clear = "none";
defparam ram_block3a32.port_b_address_clock = "clock1";
defparam ram_block3a32.port_b_address_width = 13;
defparam ram_block3a32.port_b_data_in_clock = "clock1";
defparam ram_block3a32.port_b_data_out_clear = "none";
defparam ram_block3a32.port_b_data_out_clock = "none";
defparam ram_block3a32.port_b_data_width = 1;
defparam ram_block3a32.port_b_first_address = 0;
defparam ram_block3a32.port_b_first_bit_number = 0;
defparam ram_block3a32.port_b_last_address = 8191;
defparam ram_block3a32.port_b_logical_ram_depth = 16384;
defparam ram_block3a32.port_b_logical_ram_width = 32;
defparam ram_block3a32.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a32.port_b_read_enable_clock = "clock1";
defparam ram_block3a32.port_b_write_enable_clock = "clock1";
defparam ram_block3a32.ram_block_type = "M9K";
defparam ram_block3a32.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a32.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y28_N0
cycloneive_ram_block ram_block3a0(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[0]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[0]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a0_PORTADATAOUT_bus),
	.portbdataout(ram_block3a0_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a0.clk0_core_clock_enable = "ena0";
defparam ram_block3a0.clk1_core_clock_enable = "ena1";
defparam ram_block3a0.data_interleave_offset_in_bits = 1;
defparam ram_block3a0.data_interleave_width_in_bits = 1;
defparam ram_block3a0.init_file = "meminit.hex";
defparam ram_block3a0.init_file_layout = "port_a";
defparam ram_block3a0.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a0.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a0.operation_mode = "bidir_dual_port";
defparam ram_block3a0.port_a_address_clear = "none";
defparam ram_block3a0.port_a_address_width = 13;
defparam ram_block3a0.port_a_byte_enable_clock = "none";
defparam ram_block3a0.port_a_data_out_clear = "none";
defparam ram_block3a0.port_a_data_out_clock = "none";
defparam ram_block3a0.port_a_data_width = 1;
defparam ram_block3a0.port_a_first_address = 0;
defparam ram_block3a0.port_a_first_bit_number = 0;
defparam ram_block3a0.port_a_last_address = 8191;
defparam ram_block3a0.port_a_logical_ram_depth = 16384;
defparam ram_block3a0.port_a_logical_ram_width = 32;
defparam ram_block3a0.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_address_clear = "none";
defparam ram_block3a0.port_b_address_clock = "clock1";
defparam ram_block3a0.port_b_address_width = 13;
defparam ram_block3a0.port_b_data_in_clock = "clock1";
defparam ram_block3a0.port_b_data_out_clear = "none";
defparam ram_block3a0.port_b_data_out_clock = "none";
defparam ram_block3a0.port_b_data_width = 1;
defparam ram_block3a0.port_b_first_address = 0;
defparam ram_block3a0.port_b_first_bit_number = 0;
defparam ram_block3a0.port_b_last_address = 8191;
defparam ram_block3a0.port_b_logical_ram_depth = 16384;
defparam ram_block3a0.port_b_logical_ram_width = 32;
defparam ram_block3a0.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a0.port_b_read_enable_clock = "clock1";
defparam ram_block3a0.port_b_write_enable_clock = "clock1";
defparam ram_block3a0.ram_block_type = "M9K";
defparam ram_block3a0.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a0.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001802C7EA14A7EF95C00000000000000000000000000000A242111E008528F7260;
// synopsys translate_on

// Location: M9K_X51_Y24_N0
cycloneive_ram_block ram_block3a33(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a33_PORTADATAOUT_bus),
	.portbdataout(ram_block3a33_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a33.clk0_core_clock_enable = "ena0";
defparam ram_block3a33.clk1_core_clock_enable = "ena1";
defparam ram_block3a33.data_interleave_offset_in_bits = 1;
defparam ram_block3a33.data_interleave_width_in_bits = 1;
defparam ram_block3a33.init_file = "meminit.hex";
defparam ram_block3a33.init_file_layout = "port_a";
defparam ram_block3a33.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a33.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a33.operation_mode = "bidir_dual_port";
defparam ram_block3a33.port_a_address_clear = "none";
defparam ram_block3a33.port_a_address_width = 13;
defparam ram_block3a33.port_a_byte_enable_clock = "none";
defparam ram_block3a33.port_a_data_out_clear = "none";
defparam ram_block3a33.port_a_data_out_clock = "none";
defparam ram_block3a33.port_a_data_width = 1;
defparam ram_block3a33.port_a_first_address = 0;
defparam ram_block3a33.port_a_first_bit_number = 1;
defparam ram_block3a33.port_a_last_address = 8191;
defparam ram_block3a33.port_a_logical_ram_depth = 16384;
defparam ram_block3a33.port_a_logical_ram_width = 32;
defparam ram_block3a33.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_address_clear = "none";
defparam ram_block3a33.port_b_address_clock = "clock1";
defparam ram_block3a33.port_b_address_width = 13;
defparam ram_block3a33.port_b_data_in_clock = "clock1";
defparam ram_block3a33.port_b_data_out_clear = "none";
defparam ram_block3a33.port_b_data_out_clock = "none";
defparam ram_block3a33.port_b_data_width = 1;
defparam ram_block3a33.port_b_first_address = 0;
defparam ram_block3a33.port_b_first_bit_number = 1;
defparam ram_block3a33.port_b_last_address = 8191;
defparam ram_block3a33.port_b_logical_ram_depth = 16384;
defparam ram_block3a33.port_b_logical_ram_width = 32;
defparam ram_block3a33.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a33.port_b_read_enable_clock = "clock1";
defparam ram_block3a33.port_b_write_enable_clock = "clock1";
defparam ram_block3a33.ram_block_type = "M9K";
defparam ram_block3a33.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a33.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y25_N0
cycloneive_ram_block ram_block3a1(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[1]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[1]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a1_PORTADATAOUT_bus),
	.portbdataout(ram_block3a1_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a1.clk0_core_clock_enable = "ena0";
defparam ram_block3a1.clk1_core_clock_enable = "ena1";
defparam ram_block3a1.data_interleave_offset_in_bits = 1;
defparam ram_block3a1.data_interleave_width_in_bits = 1;
defparam ram_block3a1.init_file = "meminit.hex";
defparam ram_block3a1.init_file_layout = "port_a";
defparam ram_block3a1.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a1.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a1.operation_mode = "bidir_dual_port";
defparam ram_block3a1.port_a_address_clear = "none";
defparam ram_block3a1.port_a_address_width = 13;
defparam ram_block3a1.port_a_byte_enable_clock = "none";
defparam ram_block3a1.port_a_data_out_clear = "none";
defparam ram_block3a1.port_a_data_out_clock = "none";
defparam ram_block3a1.port_a_data_width = 1;
defparam ram_block3a1.port_a_first_address = 0;
defparam ram_block3a1.port_a_first_bit_number = 1;
defparam ram_block3a1.port_a_last_address = 8191;
defparam ram_block3a1.port_a_logical_ram_depth = 16384;
defparam ram_block3a1.port_a_logical_ram_width = 32;
defparam ram_block3a1.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_address_clear = "none";
defparam ram_block3a1.port_b_address_clock = "clock1";
defparam ram_block3a1.port_b_address_width = 13;
defparam ram_block3a1.port_b_data_in_clock = "clock1";
defparam ram_block3a1.port_b_data_out_clear = "none";
defparam ram_block3a1.port_b_data_out_clock = "none";
defparam ram_block3a1.port_b_data_width = 1;
defparam ram_block3a1.port_b_first_address = 0;
defparam ram_block3a1.port_b_first_bit_number = 1;
defparam ram_block3a1.port_b_last_address = 8191;
defparam ram_block3a1.port_b_logical_ram_depth = 16384;
defparam ram_block3a1.port_b_logical_ram_width = 32;
defparam ram_block3a1.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a1.port_b_read_enable_clock = "clock1";
defparam ram_block3a1.port_b_write_enable_clock = "clock1";
defparam ram_block3a1.ram_block_type = "M9K";
defparam ram_block3a1.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a1.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001D4AE6429116B3C8A000000000000000000000000000012242108900D12808390;
// synopsys translate_on

// Location: M9K_X37_Y23_N0
cycloneive_ram_block ram_block3a34(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a34_PORTADATAOUT_bus),
	.portbdataout(ram_block3a34_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a34.clk0_core_clock_enable = "ena0";
defparam ram_block3a34.clk1_core_clock_enable = "ena1";
defparam ram_block3a34.data_interleave_offset_in_bits = 1;
defparam ram_block3a34.data_interleave_width_in_bits = 1;
defparam ram_block3a34.init_file = "meminit.hex";
defparam ram_block3a34.init_file_layout = "port_a";
defparam ram_block3a34.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a34.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a34.operation_mode = "bidir_dual_port";
defparam ram_block3a34.port_a_address_clear = "none";
defparam ram_block3a34.port_a_address_width = 13;
defparam ram_block3a34.port_a_byte_enable_clock = "none";
defparam ram_block3a34.port_a_data_out_clear = "none";
defparam ram_block3a34.port_a_data_out_clock = "none";
defparam ram_block3a34.port_a_data_width = 1;
defparam ram_block3a34.port_a_first_address = 0;
defparam ram_block3a34.port_a_first_bit_number = 2;
defparam ram_block3a34.port_a_last_address = 8191;
defparam ram_block3a34.port_a_logical_ram_depth = 16384;
defparam ram_block3a34.port_a_logical_ram_width = 32;
defparam ram_block3a34.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_address_clear = "none";
defparam ram_block3a34.port_b_address_clock = "clock1";
defparam ram_block3a34.port_b_address_width = 13;
defparam ram_block3a34.port_b_data_in_clock = "clock1";
defparam ram_block3a34.port_b_data_out_clear = "none";
defparam ram_block3a34.port_b_data_out_clock = "none";
defparam ram_block3a34.port_b_data_width = 1;
defparam ram_block3a34.port_b_first_address = 0;
defparam ram_block3a34.port_b_first_bit_number = 2;
defparam ram_block3a34.port_b_last_address = 8191;
defparam ram_block3a34.port_b_logical_ram_depth = 16384;
defparam ram_block3a34.port_b_logical_ram_width = 32;
defparam ram_block3a34.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a34.port_b_read_enable_clock = "clock1";
defparam ram_block3a34.port_b_write_enable_clock = "clock1";
defparam ram_block3a34.ram_block_type = "M9K";
defparam ram_block3a34.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a34.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y21_N0
cycloneive_ram_block ram_block3a2(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[2]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[2]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a2_PORTADATAOUT_bus),
	.portbdataout(ram_block3a2_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a2.clk0_core_clock_enable = "ena0";
defparam ram_block3a2.clk1_core_clock_enable = "ena1";
defparam ram_block3a2.data_interleave_offset_in_bits = 1;
defparam ram_block3a2.data_interleave_width_in_bits = 1;
defparam ram_block3a2.init_file = "meminit.hex";
defparam ram_block3a2.init_file_layout = "port_a";
defparam ram_block3a2.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a2.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a2.operation_mode = "bidir_dual_port";
defparam ram_block3a2.port_a_address_clear = "none";
defparam ram_block3a2.port_a_address_width = 13;
defparam ram_block3a2.port_a_byte_enable_clock = "none";
defparam ram_block3a2.port_a_data_out_clear = "none";
defparam ram_block3a2.port_a_data_out_clock = "none";
defparam ram_block3a2.port_a_data_width = 1;
defparam ram_block3a2.port_a_first_address = 0;
defparam ram_block3a2.port_a_first_bit_number = 2;
defparam ram_block3a2.port_a_last_address = 8191;
defparam ram_block3a2.port_a_logical_ram_depth = 16384;
defparam ram_block3a2.port_a_logical_ram_width = 32;
defparam ram_block3a2.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_address_clear = "none";
defparam ram_block3a2.port_b_address_clock = "clock1";
defparam ram_block3a2.port_b_address_width = 13;
defparam ram_block3a2.port_b_data_in_clock = "clock1";
defparam ram_block3a2.port_b_data_out_clear = "none";
defparam ram_block3a2.port_b_data_out_clock = "none";
defparam ram_block3a2.port_b_data_width = 1;
defparam ram_block3a2.port_b_first_address = 0;
defparam ram_block3a2.port_b_first_bit_number = 2;
defparam ram_block3a2.port_b_last_address = 8191;
defparam ram_block3a2.port_b_logical_ram_depth = 16384;
defparam ram_block3a2.port_b_logical_ram_width = 32;
defparam ram_block3a2.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a2.port_b_read_enable_clock = "clock1";
defparam ram_block3a2.port_b_write_enable_clock = "clock1";
defparam ram_block3a2.ram_block_type = "M9K";
defparam ram_block3a2.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a2.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000961CA470728D97800000000000000000000000000000172E7BD1C323272F6867;
// synopsys translate_on

// Location: M9K_X51_Y22_N0
cycloneive_ram_block ram_block3a35(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a35_PORTADATAOUT_bus),
	.portbdataout(ram_block3a35_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a35.clk0_core_clock_enable = "ena0";
defparam ram_block3a35.clk1_core_clock_enable = "ena1";
defparam ram_block3a35.data_interleave_offset_in_bits = 1;
defparam ram_block3a35.data_interleave_width_in_bits = 1;
defparam ram_block3a35.init_file = "meminit.hex";
defparam ram_block3a35.init_file_layout = "port_a";
defparam ram_block3a35.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a35.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a35.operation_mode = "bidir_dual_port";
defparam ram_block3a35.port_a_address_clear = "none";
defparam ram_block3a35.port_a_address_width = 13;
defparam ram_block3a35.port_a_byte_enable_clock = "none";
defparam ram_block3a35.port_a_data_out_clear = "none";
defparam ram_block3a35.port_a_data_out_clock = "none";
defparam ram_block3a35.port_a_data_width = 1;
defparam ram_block3a35.port_a_first_address = 0;
defparam ram_block3a35.port_a_first_bit_number = 3;
defparam ram_block3a35.port_a_last_address = 8191;
defparam ram_block3a35.port_a_logical_ram_depth = 16384;
defparam ram_block3a35.port_a_logical_ram_width = 32;
defparam ram_block3a35.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_address_clear = "none";
defparam ram_block3a35.port_b_address_clock = "clock1";
defparam ram_block3a35.port_b_address_width = 13;
defparam ram_block3a35.port_b_data_in_clock = "clock1";
defparam ram_block3a35.port_b_data_out_clear = "none";
defparam ram_block3a35.port_b_data_out_clock = "none";
defparam ram_block3a35.port_b_data_width = 1;
defparam ram_block3a35.port_b_first_address = 0;
defparam ram_block3a35.port_b_first_bit_number = 3;
defparam ram_block3a35.port_b_last_address = 8191;
defparam ram_block3a35.port_b_logical_ram_depth = 16384;
defparam ram_block3a35.port_b_logical_ram_width = 32;
defparam ram_block3a35.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a35.port_b_read_enable_clock = "clock1";
defparam ram_block3a35.port_b_write_enable_clock = "clock1";
defparam ram_block3a35.ram_block_type = "M9K";
defparam ram_block3a35.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a35.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y21_N0
cycloneive_ram_block ram_block3a3(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[3]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[3]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a3_PORTADATAOUT_bus),
	.portbdataout(ram_block3a3_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a3.clk0_core_clock_enable = "ena0";
defparam ram_block3a3.clk1_core_clock_enable = "ena1";
defparam ram_block3a3.data_interleave_offset_in_bits = 1;
defparam ram_block3a3.data_interleave_width_in_bits = 1;
defparam ram_block3a3.init_file = "meminit.hex";
defparam ram_block3a3.init_file_layout = "port_a";
defparam ram_block3a3.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a3.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a3.operation_mode = "bidir_dual_port";
defparam ram_block3a3.port_a_address_clear = "none";
defparam ram_block3a3.port_a_address_width = 13;
defparam ram_block3a3.port_a_byte_enable_clock = "none";
defparam ram_block3a3.port_a_data_out_clear = "none";
defparam ram_block3a3.port_a_data_out_clock = "none";
defparam ram_block3a3.port_a_data_width = 1;
defparam ram_block3a3.port_a_first_address = 0;
defparam ram_block3a3.port_a_first_bit_number = 3;
defparam ram_block3a3.port_a_last_address = 8191;
defparam ram_block3a3.port_a_logical_ram_depth = 16384;
defparam ram_block3a3.port_a_logical_ram_width = 32;
defparam ram_block3a3.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_address_clear = "none";
defparam ram_block3a3.port_b_address_clock = "clock1";
defparam ram_block3a3.port_b_address_width = 13;
defparam ram_block3a3.port_b_data_in_clock = "clock1";
defparam ram_block3a3.port_b_data_out_clear = "none";
defparam ram_block3a3.port_b_data_out_clock = "none";
defparam ram_block3a3.port_b_data_width = 1;
defparam ram_block3a3.port_b_first_address = 0;
defparam ram_block3a3.port_b_first_bit_number = 3;
defparam ram_block3a3.port_b_last_address = 8191;
defparam ram_block3a3.port_b_logical_ram_depth = 16384;
defparam ram_block3a3.port_b_logical_ram_width = 32;
defparam ram_block3a3.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a3.port_b_read_enable_clock = "clock1";
defparam ram_block3a3.port_b_write_enable_clock = "clock1";
defparam ram_block3a3.ram_block_type = "M9K";
defparam ram_block3a3.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a3.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000009F20E64C2468E52000000000000000000000000000022346308C62632A08083;
// synopsys translate_on

// Location: M9K_X37_Y26_N0
cycloneive_ram_block ram_block3a36(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a36_PORTADATAOUT_bus),
	.portbdataout(ram_block3a36_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a36.clk0_core_clock_enable = "ena0";
defparam ram_block3a36.clk1_core_clock_enable = "ena1";
defparam ram_block3a36.data_interleave_offset_in_bits = 1;
defparam ram_block3a36.data_interleave_width_in_bits = 1;
defparam ram_block3a36.init_file = "meminit.hex";
defparam ram_block3a36.init_file_layout = "port_a";
defparam ram_block3a36.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a36.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a36.operation_mode = "bidir_dual_port";
defparam ram_block3a36.port_a_address_clear = "none";
defparam ram_block3a36.port_a_address_width = 13;
defparam ram_block3a36.port_a_byte_enable_clock = "none";
defparam ram_block3a36.port_a_data_out_clear = "none";
defparam ram_block3a36.port_a_data_out_clock = "none";
defparam ram_block3a36.port_a_data_width = 1;
defparam ram_block3a36.port_a_first_address = 0;
defparam ram_block3a36.port_a_first_bit_number = 4;
defparam ram_block3a36.port_a_last_address = 8191;
defparam ram_block3a36.port_a_logical_ram_depth = 16384;
defparam ram_block3a36.port_a_logical_ram_width = 32;
defparam ram_block3a36.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_address_clear = "none";
defparam ram_block3a36.port_b_address_clock = "clock1";
defparam ram_block3a36.port_b_address_width = 13;
defparam ram_block3a36.port_b_data_in_clock = "clock1";
defparam ram_block3a36.port_b_data_out_clear = "none";
defparam ram_block3a36.port_b_data_out_clock = "none";
defparam ram_block3a36.port_b_data_width = 1;
defparam ram_block3a36.port_b_first_address = 0;
defparam ram_block3a36.port_b_first_bit_number = 4;
defparam ram_block3a36.port_b_last_address = 8191;
defparam ram_block3a36.port_b_logical_ram_depth = 16384;
defparam ram_block3a36.port_b_logical_ram_width = 32;
defparam ram_block3a36.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a36.port_b_read_enable_clock = "clock1";
defparam ram_block3a36.port_b_write_enable_clock = "clock1";
defparam ram_block3a36.ram_block_type = "M9K";
defparam ram_block3a36.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a36.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y27_N0
cycloneive_ram_block ram_block3a4(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[4]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[4]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a4_PORTADATAOUT_bus),
	.portbdataout(ram_block3a4_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a4.clk0_core_clock_enable = "ena0";
defparam ram_block3a4.clk1_core_clock_enable = "ena1";
defparam ram_block3a4.data_interleave_offset_in_bits = 1;
defparam ram_block3a4.data_interleave_width_in_bits = 1;
defparam ram_block3a4.init_file = "meminit.hex";
defparam ram_block3a4.init_file_layout = "port_a";
defparam ram_block3a4.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a4.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a4.operation_mode = "bidir_dual_port";
defparam ram_block3a4.port_a_address_clear = "none";
defparam ram_block3a4.port_a_address_width = 13;
defparam ram_block3a4.port_a_byte_enable_clock = "none";
defparam ram_block3a4.port_a_data_out_clear = "none";
defparam ram_block3a4.port_a_data_out_clock = "none";
defparam ram_block3a4.port_a_data_width = 1;
defparam ram_block3a4.port_a_first_address = 0;
defparam ram_block3a4.port_a_first_bit_number = 4;
defparam ram_block3a4.port_a_last_address = 8191;
defparam ram_block3a4.port_a_logical_ram_depth = 16384;
defparam ram_block3a4.port_a_logical_ram_width = 32;
defparam ram_block3a4.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_address_clear = "none";
defparam ram_block3a4.port_b_address_clock = "clock1";
defparam ram_block3a4.port_b_address_width = 13;
defparam ram_block3a4.port_b_data_in_clock = "clock1";
defparam ram_block3a4.port_b_data_out_clear = "none";
defparam ram_block3a4.port_b_data_out_clock = "none";
defparam ram_block3a4.port_b_data_width = 1;
defparam ram_block3a4.port_b_first_address = 0;
defparam ram_block3a4.port_b_first_bit_number = 4;
defparam ram_block3a4.port_b_last_address = 8191;
defparam ram_block3a4.port_b_logical_ram_depth = 16384;
defparam ram_block3a4.port_b_logical_ram_width = 32;
defparam ram_block3a4.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a4.port_b_read_enable_clock = "clock1";
defparam ram_block3a4.port_b_write_enable_clock = "clock1";
defparam ram_block3a4.ram_block_type = "M9K";
defparam ram_block3a4.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a4.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060B81842D24565BE000000000000000000000000000002242101022202208083;
// synopsys translate_on

// Location: M9K_X78_Y27_N0
cycloneive_ram_block ram_block3a37(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a37_PORTADATAOUT_bus),
	.portbdataout(ram_block3a37_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a37.clk0_core_clock_enable = "ena0";
defparam ram_block3a37.clk1_core_clock_enable = "ena1";
defparam ram_block3a37.data_interleave_offset_in_bits = 1;
defparam ram_block3a37.data_interleave_width_in_bits = 1;
defparam ram_block3a37.init_file = "meminit.hex";
defparam ram_block3a37.init_file_layout = "port_a";
defparam ram_block3a37.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a37.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a37.operation_mode = "bidir_dual_port";
defparam ram_block3a37.port_a_address_clear = "none";
defparam ram_block3a37.port_a_address_width = 13;
defparam ram_block3a37.port_a_byte_enable_clock = "none";
defparam ram_block3a37.port_a_data_out_clear = "none";
defparam ram_block3a37.port_a_data_out_clock = "none";
defparam ram_block3a37.port_a_data_width = 1;
defparam ram_block3a37.port_a_first_address = 0;
defparam ram_block3a37.port_a_first_bit_number = 5;
defparam ram_block3a37.port_a_last_address = 8191;
defparam ram_block3a37.port_a_logical_ram_depth = 16384;
defparam ram_block3a37.port_a_logical_ram_width = 32;
defparam ram_block3a37.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_address_clear = "none";
defparam ram_block3a37.port_b_address_clock = "clock1";
defparam ram_block3a37.port_b_address_width = 13;
defparam ram_block3a37.port_b_data_in_clock = "clock1";
defparam ram_block3a37.port_b_data_out_clear = "none";
defparam ram_block3a37.port_b_data_out_clock = "none";
defparam ram_block3a37.port_b_data_width = 1;
defparam ram_block3a37.port_b_first_address = 0;
defparam ram_block3a37.port_b_first_bit_number = 5;
defparam ram_block3a37.port_b_last_address = 8191;
defparam ram_block3a37.port_b_logical_ram_depth = 16384;
defparam ram_block3a37.port_b_logical_ram_width = 32;
defparam ram_block3a37.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a37.port_b_read_enable_clock = "clock1";
defparam ram_block3a37.port_b_write_enable_clock = "clock1";
defparam ram_block3a37.ram_block_type = "M9K";
defparam ram_block3a37.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a37.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y26_N0
cycloneive_ram_block ram_block3a5(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[5]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[5]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a5_PORTADATAOUT_bus),
	.portbdataout(ram_block3a5_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a5.clk0_core_clock_enable = "ena0";
defparam ram_block3a5.clk1_core_clock_enable = "ena1";
defparam ram_block3a5.data_interleave_offset_in_bits = 1;
defparam ram_block3a5.data_interleave_width_in_bits = 1;
defparam ram_block3a5.init_file = "meminit.hex";
defparam ram_block3a5.init_file_layout = "port_a";
defparam ram_block3a5.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a5.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a5.operation_mode = "bidir_dual_port";
defparam ram_block3a5.port_a_address_clear = "none";
defparam ram_block3a5.port_a_address_width = 13;
defparam ram_block3a5.port_a_byte_enable_clock = "none";
defparam ram_block3a5.port_a_data_out_clear = "none";
defparam ram_block3a5.port_a_data_out_clock = "none";
defparam ram_block3a5.port_a_data_width = 1;
defparam ram_block3a5.port_a_first_address = 0;
defparam ram_block3a5.port_a_first_bit_number = 5;
defparam ram_block3a5.port_a_last_address = 8191;
defparam ram_block3a5.port_a_logical_ram_depth = 16384;
defparam ram_block3a5.port_a_logical_ram_width = 32;
defparam ram_block3a5.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_address_clear = "none";
defparam ram_block3a5.port_b_address_clock = "clock1";
defparam ram_block3a5.port_b_address_width = 13;
defparam ram_block3a5.port_b_data_in_clock = "clock1";
defparam ram_block3a5.port_b_data_out_clear = "none";
defparam ram_block3a5.port_b_data_out_clock = "none";
defparam ram_block3a5.port_b_data_width = 1;
defparam ram_block3a5.port_b_first_address = 0;
defparam ram_block3a5.port_b_first_bit_number = 5;
defparam ram_block3a5.port_b_last_address = 8191;
defparam ram_block3a5.port_b_logical_ram_depth = 16384;
defparam ram_block3a5.port_b_logical_ram_width = 32;
defparam ram_block3a5.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a5.port_b_read_enable_clock = "clock1";
defparam ram_block3a5.port_b_write_enable_clock = "clock1";
defparam ram_block3a5.ram_block_type = "M9K";
defparam ram_block3a5.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a5.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000056414512D6B00448000000000000000000000000000002246308006652AF7263;
// synopsys translate_on

// Location: M9K_X78_Y25_N0
cycloneive_ram_block ram_block3a38(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a38_PORTADATAOUT_bus),
	.portbdataout(ram_block3a38_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a38.clk0_core_clock_enable = "ena0";
defparam ram_block3a38.clk1_core_clock_enable = "ena1";
defparam ram_block3a38.data_interleave_offset_in_bits = 1;
defparam ram_block3a38.data_interleave_width_in_bits = 1;
defparam ram_block3a38.init_file = "meminit.hex";
defparam ram_block3a38.init_file_layout = "port_a";
defparam ram_block3a38.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a38.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a38.operation_mode = "bidir_dual_port";
defparam ram_block3a38.port_a_address_clear = "none";
defparam ram_block3a38.port_a_address_width = 13;
defparam ram_block3a38.port_a_byte_enable_clock = "none";
defparam ram_block3a38.port_a_data_out_clear = "none";
defparam ram_block3a38.port_a_data_out_clock = "none";
defparam ram_block3a38.port_a_data_width = 1;
defparam ram_block3a38.port_a_first_address = 0;
defparam ram_block3a38.port_a_first_bit_number = 6;
defparam ram_block3a38.port_a_last_address = 8191;
defparam ram_block3a38.port_a_logical_ram_depth = 16384;
defparam ram_block3a38.port_a_logical_ram_width = 32;
defparam ram_block3a38.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_address_clear = "none";
defparam ram_block3a38.port_b_address_clock = "clock1";
defparam ram_block3a38.port_b_address_width = 13;
defparam ram_block3a38.port_b_data_in_clock = "clock1";
defparam ram_block3a38.port_b_data_out_clear = "none";
defparam ram_block3a38.port_b_data_out_clock = "none";
defparam ram_block3a38.port_b_data_width = 1;
defparam ram_block3a38.port_b_first_address = 0;
defparam ram_block3a38.port_b_first_bit_number = 6;
defparam ram_block3a38.port_b_last_address = 8191;
defparam ram_block3a38.port_b_logical_ram_depth = 16384;
defparam ram_block3a38.port_b_logical_ram_width = 32;
defparam ram_block3a38.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a38.port_b_read_enable_clock = "clock1";
defparam ram_block3a38.port_b_write_enable_clock = "clock1";
defparam ram_block3a38.ram_block_type = "M9K";
defparam ram_block3a38.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a38.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y28_N0
cycloneive_ram_block ram_block3a6(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[6]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[6]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a6_PORTADATAOUT_bus),
	.portbdataout(ram_block3a6_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a6.clk0_core_clock_enable = "ena0";
defparam ram_block3a6.clk1_core_clock_enable = "ena1";
defparam ram_block3a6.data_interleave_offset_in_bits = 1;
defparam ram_block3a6.data_interleave_width_in_bits = 1;
defparam ram_block3a6.init_file = "meminit.hex";
defparam ram_block3a6.init_file_layout = "port_a";
defparam ram_block3a6.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a6.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a6.operation_mode = "bidir_dual_port";
defparam ram_block3a6.port_a_address_clear = "none";
defparam ram_block3a6.port_a_address_width = 13;
defparam ram_block3a6.port_a_byte_enable_clock = "none";
defparam ram_block3a6.port_a_data_out_clear = "none";
defparam ram_block3a6.port_a_data_out_clock = "none";
defparam ram_block3a6.port_a_data_width = 1;
defparam ram_block3a6.port_a_first_address = 0;
defparam ram_block3a6.port_a_first_bit_number = 6;
defparam ram_block3a6.port_a_last_address = 8191;
defparam ram_block3a6.port_a_logical_ram_depth = 16384;
defparam ram_block3a6.port_a_logical_ram_width = 32;
defparam ram_block3a6.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_address_clear = "none";
defparam ram_block3a6.port_b_address_clock = "clock1";
defparam ram_block3a6.port_b_address_width = 13;
defparam ram_block3a6.port_b_data_in_clock = "clock1";
defparam ram_block3a6.port_b_data_out_clear = "none";
defparam ram_block3a6.port_b_data_out_clock = "none";
defparam ram_block3a6.port_b_data_width = 1;
defparam ram_block3a6.port_b_first_address = 0;
defparam ram_block3a6.port_b_first_bit_number = 6;
defparam ram_block3a6.port_b_last_address = 8191;
defparam ram_block3a6.port_b_logical_ram_depth = 16384;
defparam ram_block3a6.port_b_logical_ram_width = 32;
defparam ram_block3a6.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a6.port_b_read_enable_clock = "clock1";
defparam ram_block3a6.port_b_write_enable_clock = "clock1";
defparam ram_block3a6.ram_block_type = "M9K";
defparam ram_block3a6.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a6.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001003088D801A0F827000000000000000000000000000012042100402202200113;
// synopsys translate_on

// Location: M9K_X64_Y23_N0
cycloneive_ram_block ram_block3a39(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a39_PORTADATAOUT_bus),
	.portbdataout(ram_block3a39_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a39.clk0_core_clock_enable = "ena0";
defparam ram_block3a39.clk1_core_clock_enable = "ena1";
defparam ram_block3a39.data_interleave_offset_in_bits = 1;
defparam ram_block3a39.data_interleave_width_in_bits = 1;
defparam ram_block3a39.init_file = "meminit.hex";
defparam ram_block3a39.init_file_layout = "port_a";
defparam ram_block3a39.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a39.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a39.operation_mode = "bidir_dual_port";
defparam ram_block3a39.port_a_address_clear = "none";
defparam ram_block3a39.port_a_address_width = 13;
defparam ram_block3a39.port_a_byte_enable_clock = "none";
defparam ram_block3a39.port_a_data_out_clear = "none";
defparam ram_block3a39.port_a_data_out_clock = "none";
defparam ram_block3a39.port_a_data_width = 1;
defparam ram_block3a39.port_a_first_address = 0;
defparam ram_block3a39.port_a_first_bit_number = 7;
defparam ram_block3a39.port_a_last_address = 8191;
defparam ram_block3a39.port_a_logical_ram_depth = 16384;
defparam ram_block3a39.port_a_logical_ram_width = 32;
defparam ram_block3a39.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_address_clear = "none";
defparam ram_block3a39.port_b_address_clock = "clock1";
defparam ram_block3a39.port_b_address_width = 13;
defparam ram_block3a39.port_b_data_in_clock = "clock1";
defparam ram_block3a39.port_b_data_out_clear = "none";
defparam ram_block3a39.port_b_data_out_clock = "none";
defparam ram_block3a39.port_b_data_width = 1;
defparam ram_block3a39.port_b_first_address = 0;
defparam ram_block3a39.port_b_first_bit_number = 7;
defparam ram_block3a39.port_b_last_address = 8191;
defparam ram_block3a39.port_b_logical_ram_depth = 16384;
defparam ram_block3a39.port_b_logical_ram_width = 32;
defparam ram_block3a39.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a39.port_b_read_enable_clock = "clock1";
defparam ram_block3a39.port_b_write_enable_clock = "clock1";
defparam ram_block3a39.ram_block_type = "M9K";
defparam ram_block3a39.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a39.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y23_N0
cycloneive_ram_block ram_block3a7(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[7]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[7]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a7_PORTADATAOUT_bus),
	.portbdataout(ram_block3a7_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a7.clk0_core_clock_enable = "ena0";
defparam ram_block3a7.clk1_core_clock_enable = "ena1";
defparam ram_block3a7.data_interleave_offset_in_bits = 1;
defparam ram_block3a7.data_interleave_width_in_bits = 1;
defparam ram_block3a7.init_file = "meminit.hex";
defparam ram_block3a7.init_file_layout = "port_a";
defparam ram_block3a7.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a7.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a7.operation_mode = "bidir_dual_port";
defparam ram_block3a7.port_a_address_clear = "none";
defparam ram_block3a7.port_a_address_width = 13;
defparam ram_block3a7.port_a_byte_enable_clock = "none";
defparam ram_block3a7.port_a_data_out_clear = "none";
defparam ram_block3a7.port_a_data_out_clock = "none";
defparam ram_block3a7.port_a_data_width = 1;
defparam ram_block3a7.port_a_first_address = 0;
defparam ram_block3a7.port_a_first_bit_number = 7;
defparam ram_block3a7.port_a_last_address = 8191;
defparam ram_block3a7.port_a_logical_ram_depth = 16384;
defparam ram_block3a7.port_a_logical_ram_width = 32;
defparam ram_block3a7.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_address_clear = "none";
defparam ram_block3a7.port_b_address_clock = "clock1";
defparam ram_block3a7.port_b_address_width = 13;
defparam ram_block3a7.port_b_data_in_clock = "clock1";
defparam ram_block3a7.port_b_data_out_clear = "none";
defparam ram_block3a7.port_b_data_out_clock = "none";
defparam ram_block3a7.port_b_data_width = 1;
defparam ram_block3a7.port_b_first_address = 0;
defparam ram_block3a7.port_b_first_bit_number = 7;
defparam ram_block3a7.port_b_last_address = 8191;
defparam ram_block3a7.port_b_logical_ram_depth = 16384;
defparam ram_block3a7.port_b_logical_ram_width = 32;
defparam ram_block3a7.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a7.port_b_read_enable_clock = "clock1";
defparam ram_block3a7.port_b_write_enable_clock = "clock1";
defparam ram_block3a7.ram_block_type = "M9K";
defparam ram_block3a7.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a7.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220A200403;
// synopsys translate_on

// Location: M9K_X64_Y27_N0
cycloneive_ram_block ram_block3a40(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a40_PORTADATAOUT_bus),
	.portbdataout(ram_block3a40_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a40.clk0_core_clock_enable = "ena0";
defparam ram_block3a40.clk1_core_clock_enable = "ena1";
defparam ram_block3a40.data_interleave_offset_in_bits = 1;
defparam ram_block3a40.data_interleave_width_in_bits = 1;
defparam ram_block3a40.init_file = "meminit.hex";
defparam ram_block3a40.init_file_layout = "port_a";
defparam ram_block3a40.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a40.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a40.operation_mode = "bidir_dual_port";
defparam ram_block3a40.port_a_address_clear = "none";
defparam ram_block3a40.port_a_address_width = 13;
defparam ram_block3a40.port_a_byte_enable_clock = "none";
defparam ram_block3a40.port_a_data_out_clear = "none";
defparam ram_block3a40.port_a_data_out_clock = "none";
defparam ram_block3a40.port_a_data_width = 1;
defparam ram_block3a40.port_a_first_address = 0;
defparam ram_block3a40.port_a_first_bit_number = 8;
defparam ram_block3a40.port_a_last_address = 8191;
defparam ram_block3a40.port_a_logical_ram_depth = 16384;
defparam ram_block3a40.port_a_logical_ram_width = 32;
defparam ram_block3a40.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_address_clear = "none";
defparam ram_block3a40.port_b_address_clock = "clock1";
defparam ram_block3a40.port_b_address_width = 13;
defparam ram_block3a40.port_b_data_in_clock = "clock1";
defparam ram_block3a40.port_b_data_out_clear = "none";
defparam ram_block3a40.port_b_data_out_clock = "none";
defparam ram_block3a40.port_b_data_width = 1;
defparam ram_block3a40.port_b_first_address = 0;
defparam ram_block3a40.port_b_first_bit_number = 8;
defparam ram_block3a40.port_b_last_address = 8191;
defparam ram_block3a40.port_b_logical_ram_depth = 16384;
defparam ram_block3a40.port_b_logical_ram_width = 32;
defparam ram_block3a40.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a40.port_b_read_enable_clock = "clock1";
defparam ram_block3a40.port_b_write_enable_clock = "clock1";
defparam ram_block3a40.ram_block_type = "M9K";
defparam ram_block3a40.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a40.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y26_N0
cycloneive_ram_block ram_block3a8(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[8]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[8]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a8_PORTADATAOUT_bus),
	.portbdataout(ram_block3a8_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a8.clk0_core_clock_enable = "ena0";
defparam ram_block3a8.clk1_core_clock_enable = "ena1";
defparam ram_block3a8.data_interleave_offset_in_bits = 1;
defparam ram_block3a8.data_interleave_width_in_bits = 1;
defparam ram_block3a8.init_file = "meminit.hex";
defparam ram_block3a8.init_file_layout = "port_a";
defparam ram_block3a8.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a8.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a8.operation_mode = "bidir_dual_port";
defparam ram_block3a8.port_a_address_clear = "none";
defparam ram_block3a8.port_a_address_width = 13;
defparam ram_block3a8.port_a_byte_enable_clock = "none";
defparam ram_block3a8.port_a_data_out_clear = "none";
defparam ram_block3a8.port_a_data_out_clock = "none";
defparam ram_block3a8.port_a_data_width = 1;
defparam ram_block3a8.port_a_first_address = 0;
defparam ram_block3a8.port_a_first_bit_number = 8;
defparam ram_block3a8.port_a_last_address = 8191;
defparam ram_block3a8.port_a_logical_ram_depth = 16384;
defparam ram_block3a8.port_a_logical_ram_width = 32;
defparam ram_block3a8.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_address_clear = "none";
defparam ram_block3a8.port_b_address_clock = "clock1";
defparam ram_block3a8.port_b_address_width = 13;
defparam ram_block3a8.port_b_data_in_clock = "clock1";
defparam ram_block3a8.port_b_data_out_clear = "none";
defparam ram_block3a8.port_b_data_out_clock = "none";
defparam ram_block3a8.port_b_data_width = 1;
defparam ram_block3a8.port_b_first_address = 0;
defparam ram_block3a8.port_b_first_bit_number = 8;
defparam ram_block3a8.port_b_last_address = 8191;
defparam ram_block3a8.port_b_logical_ram_depth = 16384;
defparam ram_block3a8.port_b_logical_ram_width = 32;
defparam ram_block3a8.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a8.port_b_read_enable_clock = "clock1";
defparam ram_block3a8.port_b_write_enable_clock = "clock1";
defparam ram_block3a8.ram_block_type = "M9K";
defparam ram_block3a8.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a8.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220230080F;
// synopsys translate_on

// Location: M9K_X37_Y25_N0
cycloneive_ram_block ram_block3a41(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a41_PORTADATAOUT_bus),
	.portbdataout(ram_block3a41_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a41.clk0_core_clock_enable = "ena0";
defparam ram_block3a41.clk1_core_clock_enable = "ena1";
defparam ram_block3a41.data_interleave_offset_in_bits = 1;
defparam ram_block3a41.data_interleave_width_in_bits = 1;
defparam ram_block3a41.init_file = "meminit.hex";
defparam ram_block3a41.init_file_layout = "port_a";
defparam ram_block3a41.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a41.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a41.operation_mode = "bidir_dual_port";
defparam ram_block3a41.port_a_address_clear = "none";
defparam ram_block3a41.port_a_address_width = 13;
defparam ram_block3a41.port_a_byte_enable_clock = "none";
defparam ram_block3a41.port_a_data_out_clear = "none";
defparam ram_block3a41.port_a_data_out_clock = "none";
defparam ram_block3a41.port_a_data_width = 1;
defparam ram_block3a41.port_a_first_address = 0;
defparam ram_block3a41.port_a_first_bit_number = 9;
defparam ram_block3a41.port_a_last_address = 8191;
defparam ram_block3a41.port_a_logical_ram_depth = 16384;
defparam ram_block3a41.port_a_logical_ram_width = 32;
defparam ram_block3a41.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_address_clear = "none";
defparam ram_block3a41.port_b_address_clock = "clock1";
defparam ram_block3a41.port_b_address_width = 13;
defparam ram_block3a41.port_b_data_in_clock = "clock1";
defparam ram_block3a41.port_b_data_out_clear = "none";
defparam ram_block3a41.port_b_data_out_clock = "none";
defparam ram_block3a41.port_b_data_width = 1;
defparam ram_block3a41.port_b_first_address = 0;
defparam ram_block3a41.port_b_first_bit_number = 9;
defparam ram_block3a41.port_b_last_address = 8191;
defparam ram_block3a41.port_b_logical_ram_depth = 16384;
defparam ram_block3a41.port_b_logical_ram_width = 32;
defparam ram_block3a41.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a41.port_b_read_enable_clock = "clock1";
defparam ram_block3a41.port_b_write_enable_clock = "clock1";
defparam ram_block3a41.ram_block_type = "M9K";
defparam ram_block3a41.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a41.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y24_N0
cycloneive_ram_block ram_block3a9(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[9]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[9]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a9_PORTADATAOUT_bus),
	.portbdataout(ram_block3a9_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a9.clk0_core_clock_enable = "ena0";
defparam ram_block3a9.clk1_core_clock_enable = "ena1";
defparam ram_block3a9.data_interleave_offset_in_bits = 1;
defparam ram_block3a9.data_interleave_width_in_bits = 1;
defparam ram_block3a9.init_file = "meminit.hex";
defparam ram_block3a9.init_file_layout = "port_a";
defparam ram_block3a9.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a9.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a9.operation_mode = "bidir_dual_port";
defparam ram_block3a9.port_a_address_clear = "none";
defparam ram_block3a9.port_a_address_width = 13;
defparam ram_block3a9.port_a_byte_enable_clock = "none";
defparam ram_block3a9.port_a_data_out_clear = "none";
defparam ram_block3a9.port_a_data_out_clock = "none";
defparam ram_block3a9.port_a_data_width = 1;
defparam ram_block3a9.port_a_first_address = 0;
defparam ram_block3a9.port_a_first_bit_number = 9;
defparam ram_block3a9.port_a_last_address = 8191;
defparam ram_block3a9.port_a_logical_ram_depth = 16384;
defparam ram_block3a9.port_a_logical_ram_width = 32;
defparam ram_block3a9.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_address_clear = "none";
defparam ram_block3a9.port_b_address_clock = "clock1";
defparam ram_block3a9.port_b_address_width = 13;
defparam ram_block3a9.port_b_data_in_clock = "clock1";
defparam ram_block3a9.port_b_data_out_clear = "none";
defparam ram_block3a9.port_b_data_out_clock = "none";
defparam ram_block3a9.port_b_data_width = 1;
defparam ram_block3a9.port_b_first_address = 0;
defparam ram_block3a9.port_b_first_bit_number = 9;
defparam ram_block3a9.port_b_last_address = 8191;
defparam ram_block3a9.port_b_logical_ram_depth = 16384;
defparam ram_block3a9.port_b_logical_ram_width = 32;
defparam ram_block3a9.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a9.port_b_read_enable_clock = "clock1";
defparam ram_block3a9.port_b_write_enable_clock = "clock1";
defparam ram_block3a9.ram_block_type = "M9K";
defparam ram_block3a9.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a9.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000220220080F;
// synopsys translate_on

// Location: M9K_X78_Y31_N0
cycloneive_ram_block ram_block3a42(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a42_PORTADATAOUT_bus),
	.portbdataout(ram_block3a42_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a42.clk0_core_clock_enable = "ena0";
defparam ram_block3a42.clk1_core_clock_enable = "ena1";
defparam ram_block3a42.data_interleave_offset_in_bits = 1;
defparam ram_block3a42.data_interleave_width_in_bits = 1;
defparam ram_block3a42.init_file = "meminit.hex";
defparam ram_block3a42.init_file_layout = "port_a";
defparam ram_block3a42.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a42.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a42.operation_mode = "bidir_dual_port";
defparam ram_block3a42.port_a_address_clear = "none";
defparam ram_block3a42.port_a_address_width = 13;
defparam ram_block3a42.port_a_byte_enable_clock = "none";
defparam ram_block3a42.port_a_data_out_clear = "none";
defparam ram_block3a42.port_a_data_out_clock = "none";
defparam ram_block3a42.port_a_data_width = 1;
defparam ram_block3a42.port_a_first_address = 0;
defparam ram_block3a42.port_a_first_bit_number = 10;
defparam ram_block3a42.port_a_last_address = 8191;
defparam ram_block3a42.port_a_logical_ram_depth = 16384;
defparam ram_block3a42.port_a_logical_ram_width = 32;
defparam ram_block3a42.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_address_clear = "none";
defparam ram_block3a42.port_b_address_clock = "clock1";
defparam ram_block3a42.port_b_address_width = 13;
defparam ram_block3a42.port_b_data_in_clock = "clock1";
defparam ram_block3a42.port_b_data_out_clear = "none";
defparam ram_block3a42.port_b_data_out_clock = "none";
defparam ram_block3a42.port_b_data_width = 1;
defparam ram_block3a42.port_b_first_address = 0;
defparam ram_block3a42.port_b_first_bit_number = 10;
defparam ram_block3a42.port_b_last_address = 8191;
defparam ram_block3a42.port_b_logical_ram_depth = 16384;
defparam ram_block3a42.port_b_logical_ram_width = 32;
defparam ram_block3a42.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a42.port_b_read_enable_clock = "clock1";
defparam ram_block3a42.port_b_write_enable_clock = "clock1";
defparam ram_block3a42.ram_block_type = "M9K";
defparam ram_block3a42.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a42.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y34_N0
cycloneive_ram_block ram_block3a10(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[10]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[10]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a10_PORTADATAOUT_bus),
	.portbdataout(ram_block3a10_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a10.clk0_core_clock_enable = "ena0";
defparam ram_block3a10.clk1_core_clock_enable = "ena1";
defparam ram_block3a10.data_interleave_offset_in_bits = 1;
defparam ram_block3a10.data_interleave_width_in_bits = 1;
defparam ram_block3a10.init_file = "meminit.hex";
defparam ram_block3a10.init_file_layout = "port_a";
defparam ram_block3a10.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a10.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a10.operation_mode = "bidir_dual_port";
defparam ram_block3a10.port_a_address_clear = "none";
defparam ram_block3a10.port_a_address_width = 13;
defparam ram_block3a10.port_a_byte_enable_clock = "none";
defparam ram_block3a10.port_a_data_out_clear = "none";
defparam ram_block3a10.port_a_data_out_clock = "none";
defparam ram_block3a10.port_a_data_width = 1;
defparam ram_block3a10.port_a_first_address = 0;
defparam ram_block3a10.port_a_first_bit_number = 10;
defparam ram_block3a10.port_a_last_address = 8191;
defparam ram_block3a10.port_a_logical_ram_depth = 16384;
defparam ram_block3a10.port_a_logical_ram_width = 32;
defparam ram_block3a10.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_address_clear = "none";
defparam ram_block3a10.port_b_address_clock = "clock1";
defparam ram_block3a10.port_b_address_width = 13;
defparam ram_block3a10.port_b_data_in_clock = "clock1";
defparam ram_block3a10.port_b_data_out_clear = "none";
defparam ram_block3a10.port_b_data_out_clock = "none";
defparam ram_block3a10.port_b_data_width = 1;
defparam ram_block3a10.port_b_first_address = 0;
defparam ram_block3a10.port_b_first_bit_number = 10;
defparam ram_block3a10.port_b_last_address = 8191;
defparam ram_block3a10.port_b_logical_ram_depth = 16384;
defparam ram_block3a10.port_b_logical_ram_width = 32;
defparam ram_block3a10.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a10.port_b_read_enable_clock = "clock1";
defparam ram_block3a10.port_b_write_enable_clock = "clock1";
defparam ram_block3a10.ram_block_type = "M9K";
defparam ram_block3a10.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a10.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002202300003;
// synopsys translate_on

// Location: M9K_X78_Y33_N0
cycloneive_ram_block ram_block3a43(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a43_PORTADATAOUT_bus),
	.portbdataout(ram_block3a43_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a43.clk0_core_clock_enable = "ena0";
defparam ram_block3a43.clk1_core_clock_enable = "ena1";
defparam ram_block3a43.data_interleave_offset_in_bits = 1;
defparam ram_block3a43.data_interleave_width_in_bits = 1;
defparam ram_block3a43.init_file = "meminit.hex";
defparam ram_block3a43.init_file_layout = "port_a";
defparam ram_block3a43.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a43.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a43.operation_mode = "bidir_dual_port";
defparam ram_block3a43.port_a_address_clear = "none";
defparam ram_block3a43.port_a_address_width = 13;
defparam ram_block3a43.port_a_byte_enable_clock = "none";
defparam ram_block3a43.port_a_data_out_clear = "none";
defparam ram_block3a43.port_a_data_out_clock = "none";
defparam ram_block3a43.port_a_data_width = 1;
defparam ram_block3a43.port_a_first_address = 0;
defparam ram_block3a43.port_a_first_bit_number = 11;
defparam ram_block3a43.port_a_last_address = 8191;
defparam ram_block3a43.port_a_logical_ram_depth = 16384;
defparam ram_block3a43.port_a_logical_ram_width = 32;
defparam ram_block3a43.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_address_clear = "none";
defparam ram_block3a43.port_b_address_clock = "clock1";
defparam ram_block3a43.port_b_address_width = 13;
defparam ram_block3a43.port_b_data_in_clock = "clock1";
defparam ram_block3a43.port_b_data_out_clear = "none";
defparam ram_block3a43.port_b_data_out_clock = "none";
defparam ram_block3a43.port_b_data_width = 1;
defparam ram_block3a43.port_b_first_address = 0;
defparam ram_block3a43.port_b_first_bit_number = 11;
defparam ram_block3a43.port_b_last_address = 8191;
defparam ram_block3a43.port_b_logical_ram_depth = 16384;
defparam ram_block3a43.port_b_logical_ram_width = 32;
defparam ram_block3a43.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a43.port_b_read_enable_clock = "clock1";
defparam ram_block3a43.port_b_write_enable_clock = "clock1";
defparam ram_block3a43.ram_block_type = "M9K";
defparam ram_block3a43.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a43.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y35_N0
cycloneive_ram_block ram_block3a11(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[11]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[11]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a11_PORTADATAOUT_bus),
	.portbdataout(ram_block3a11_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a11.clk0_core_clock_enable = "ena0";
defparam ram_block3a11.clk1_core_clock_enable = "ena1";
defparam ram_block3a11.data_interleave_offset_in_bits = 1;
defparam ram_block3a11.data_interleave_width_in_bits = 1;
defparam ram_block3a11.init_file = "meminit.hex";
defparam ram_block3a11.init_file_layout = "port_a";
defparam ram_block3a11.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a11.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a11.operation_mode = "bidir_dual_port";
defparam ram_block3a11.port_a_address_clear = "none";
defparam ram_block3a11.port_a_address_width = 13;
defparam ram_block3a11.port_a_byte_enable_clock = "none";
defparam ram_block3a11.port_a_data_out_clear = "none";
defparam ram_block3a11.port_a_data_out_clock = "none";
defparam ram_block3a11.port_a_data_width = 1;
defparam ram_block3a11.port_a_first_address = 0;
defparam ram_block3a11.port_a_first_bit_number = 11;
defparam ram_block3a11.port_a_last_address = 8191;
defparam ram_block3a11.port_a_logical_ram_depth = 16384;
defparam ram_block3a11.port_a_logical_ram_width = 32;
defparam ram_block3a11.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_address_clear = "none";
defparam ram_block3a11.port_b_address_clock = "clock1";
defparam ram_block3a11.port_b_address_width = 13;
defparam ram_block3a11.port_b_data_in_clock = "clock1";
defparam ram_block3a11.port_b_data_out_clear = "none";
defparam ram_block3a11.port_b_data_out_clock = "none";
defparam ram_block3a11.port_b_data_width = 1;
defparam ram_block3a11.port_b_first_address = 0;
defparam ram_block3a11.port_b_first_bit_number = 11;
defparam ram_block3a11.port_b_last_address = 8191;
defparam ram_block3a11.port_b_logical_ram_depth = 16384;
defparam ram_block3a11.port_b_logical_ram_width = 32;
defparam ram_block3a11.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a11.port_b_read_enable_clock = "clock1";
defparam ram_block3a11.port_b_write_enable_clock = "clock1";
defparam ram_block3a11.ram_block_type = "M9K";
defparam ram_block3a11.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a11.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210800265A2A2233;
// synopsys translate_on

// Location: M9K_X78_Y32_N0
cycloneive_ram_block ram_block3a44(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a44_PORTADATAOUT_bus),
	.portbdataout(ram_block3a44_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a44.clk0_core_clock_enable = "ena0";
defparam ram_block3a44.clk1_core_clock_enable = "ena1";
defparam ram_block3a44.data_interleave_offset_in_bits = 1;
defparam ram_block3a44.data_interleave_width_in_bits = 1;
defparam ram_block3a44.init_file = "meminit.hex";
defparam ram_block3a44.init_file_layout = "port_a";
defparam ram_block3a44.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a44.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a44.operation_mode = "bidir_dual_port";
defparam ram_block3a44.port_a_address_clear = "none";
defparam ram_block3a44.port_a_address_width = 13;
defparam ram_block3a44.port_a_byte_enable_clock = "none";
defparam ram_block3a44.port_a_data_out_clear = "none";
defparam ram_block3a44.port_a_data_out_clock = "none";
defparam ram_block3a44.port_a_data_width = 1;
defparam ram_block3a44.port_a_first_address = 0;
defparam ram_block3a44.port_a_first_bit_number = 12;
defparam ram_block3a44.port_a_last_address = 8191;
defparam ram_block3a44.port_a_logical_ram_depth = 16384;
defparam ram_block3a44.port_a_logical_ram_width = 32;
defparam ram_block3a44.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_address_clear = "none";
defparam ram_block3a44.port_b_address_clock = "clock1";
defparam ram_block3a44.port_b_address_width = 13;
defparam ram_block3a44.port_b_data_in_clock = "clock1";
defparam ram_block3a44.port_b_data_out_clear = "none";
defparam ram_block3a44.port_b_data_out_clock = "none";
defparam ram_block3a44.port_b_data_width = 1;
defparam ram_block3a44.port_b_first_address = 0;
defparam ram_block3a44.port_b_first_bit_number = 12;
defparam ram_block3a44.port_b_last_address = 8191;
defparam ram_block3a44.port_b_logical_ram_depth = 16384;
defparam ram_block3a44.port_b_logical_ram_width = 32;
defparam ram_block3a44.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a44.port_b_read_enable_clock = "clock1";
defparam ram_block3a44.port_b_write_enable_clock = "clock1";
defparam ram_block3a44.ram_block_type = "M9K";
defparam ram_block3a44.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a44.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y29_N0
cycloneive_ram_block ram_block3a12(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[12]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[12]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a12_PORTADATAOUT_bus),
	.portbdataout(ram_block3a12_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a12.clk0_core_clock_enable = "ena0";
defparam ram_block3a12.clk1_core_clock_enable = "ena1";
defparam ram_block3a12.data_interleave_offset_in_bits = 1;
defparam ram_block3a12.data_interleave_width_in_bits = 1;
defparam ram_block3a12.init_file = "meminit.hex";
defparam ram_block3a12.init_file_layout = "port_a";
defparam ram_block3a12.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a12.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a12.operation_mode = "bidir_dual_port";
defparam ram_block3a12.port_a_address_clear = "none";
defparam ram_block3a12.port_a_address_width = 13;
defparam ram_block3a12.port_a_byte_enable_clock = "none";
defparam ram_block3a12.port_a_data_out_clear = "none";
defparam ram_block3a12.port_a_data_out_clock = "none";
defparam ram_block3a12.port_a_data_width = 1;
defparam ram_block3a12.port_a_first_address = 0;
defparam ram_block3a12.port_a_first_bit_number = 12;
defparam ram_block3a12.port_a_last_address = 8191;
defparam ram_block3a12.port_a_logical_ram_depth = 16384;
defparam ram_block3a12.port_a_logical_ram_width = 32;
defparam ram_block3a12.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_address_clear = "none";
defparam ram_block3a12.port_b_address_clock = "clock1";
defparam ram_block3a12.port_b_address_width = 13;
defparam ram_block3a12.port_b_data_in_clock = "clock1";
defparam ram_block3a12.port_b_data_out_clear = "none";
defparam ram_block3a12.port_b_data_out_clock = "none";
defparam ram_block3a12.port_b_data_width = 1;
defparam ram_block3a12.port_b_first_address = 0;
defparam ram_block3a12.port_b_first_bit_number = 12;
defparam ram_block3a12.port_b_last_address = 8191;
defparam ram_block3a12.port_b_logical_ram_depth = 16384;
defparam ram_block3a12.port_b_logical_ram_width = 32;
defparam ram_block3a12.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a12.port_b_read_enable_clock = "clock1";
defparam ram_block3a12.port_b_write_enable_clock = "clock1";
defparam ram_block3a12.ram_block_type = "M9K";
defparam ram_block3a12.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a12.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022C2043;
// synopsys translate_on

// Location: M9K_X64_Y25_N0
cycloneive_ram_block ram_block3a45(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a45_PORTADATAOUT_bus),
	.portbdataout(ram_block3a45_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a45.clk0_core_clock_enable = "ena0";
defparam ram_block3a45.clk1_core_clock_enable = "ena1";
defparam ram_block3a45.data_interleave_offset_in_bits = 1;
defparam ram_block3a45.data_interleave_width_in_bits = 1;
defparam ram_block3a45.init_file = "meminit.hex";
defparam ram_block3a45.init_file_layout = "port_a";
defparam ram_block3a45.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a45.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a45.operation_mode = "bidir_dual_port";
defparam ram_block3a45.port_a_address_clear = "none";
defparam ram_block3a45.port_a_address_width = 13;
defparam ram_block3a45.port_a_byte_enable_clock = "none";
defparam ram_block3a45.port_a_data_out_clear = "none";
defparam ram_block3a45.port_a_data_out_clock = "none";
defparam ram_block3a45.port_a_data_width = 1;
defparam ram_block3a45.port_a_first_address = 0;
defparam ram_block3a45.port_a_first_bit_number = 13;
defparam ram_block3a45.port_a_last_address = 8191;
defparam ram_block3a45.port_a_logical_ram_depth = 16384;
defparam ram_block3a45.port_a_logical_ram_width = 32;
defparam ram_block3a45.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_address_clear = "none";
defparam ram_block3a45.port_b_address_clock = "clock1";
defparam ram_block3a45.port_b_address_width = 13;
defparam ram_block3a45.port_b_data_in_clock = "clock1";
defparam ram_block3a45.port_b_data_out_clear = "none";
defparam ram_block3a45.port_b_data_out_clock = "none";
defparam ram_block3a45.port_b_data_width = 1;
defparam ram_block3a45.port_b_first_address = 0;
defparam ram_block3a45.port_b_first_bit_number = 13;
defparam ram_block3a45.port_b_last_address = 8191;
defparam ram_block3a45.port_b_logical_ram_depth = 16384;
defparam ram_block3a45.port_b_logical_ram_width = 32;
defparam ram_block3a45.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a45.port_b_read_enable_clock = "clock1";
defparam ram_block3a45.port_b_write_enable_clock = "clock1";
defparam ram_block3a45.ram_block_type = "M9K";
defparam ram_block3a45.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a45.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y26_N0
cycloneive_ram_block ram_block3a13(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[13]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[13]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a13_PORTADATAOUT_bus),
	.portbdataout(ram_block3a13_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a13.clk0_core_clock_enable = "ena0";
defparam ram_block3a13.clk1_core_clock_enable = "ena1";
defparam ram_block3a13.data_interleave_offset_in_bits = 1;
defparam ram_block3a13.data_interleave_width_in_bits = 1;
defparam ram_block3a13.init_file = "meminit.hex";
defparam ram_block3a13.init_file_layout = "port_a";
defparam ram_block3a13.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a13.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a13.operation_mode = "bidir_dual_port";
defparam ram_block3a13.port_a_address_clear = "none";
defparam ram_block3a13.port_a_address_width = 13;
defparam ram_block3a13.port_a_byte_enable_clock = "none";
defparam ram_block3a13.port_a_data_out_clear = "none";
defparam ram_block3a13.port_a_data_out_clock = "none";
defparam ram_block3a13.port_a_data_width = 1;
defparam ram_block3a13.port_a_first_address = 0;
defparam ram_block3a13.port_a_first_bit_number = 13;
defparam ram_block3a13.port_a_last_address = 8191;
defparam ram_block3a13.port_a_logical_ram_depth = 16384;
defparam ram_block3a13.port_a_logical_ram_width = 32;
defparam ram_block3a13.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_address_clear = "none";
defparam ram_block3a13.port_b_address_clock = "clock1";
defparam ram_block3a13.port_b_address_width = 13;
defparam ram_block3a13.port_b_data_in_clock = "clock1";
defparam ram_block3a13.port_b_data_out_clear = "none";
defparam ram_block3a13.port_b_data_out_clock = "none";
defparam ram_block3a13.port_b_data_width = 1;
defparam ram_block3a13.port_b_first_address = 0;
defparam ram_block3a13.port_b_first_bit_number = 13;
defparam ram_block3a13.port_b_last_address = 8191;
defparam ram_block3a13.port_b_logical_ram_depth = 16384;
defparam ram_block3a13.port_b_logical_ram_width = 32;
defparam ram_block3a13.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a13.port_b_read_enable_clock = "clock1";
defparam ram_block3a13.port_b_write_enable_clock = "clock1";
defparam ram_block3a13.ram_block_type = "M9K";
defparam ram_block3a13.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a13.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000020421000022022F5213;
// synopsys translate_on

// Location: M9K_X78_Y30_N0
cycloneive_ram_block ram_block3a46(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a46_PORTADATAOUT_bus),
	.portbdataout(ram_block3a46_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a46.clk0_core_clock_enable = "ena0";
defparam ram_block3a46.clk1_core_clock_enable = "ena1";
defparam ram_block3a46.data_interleave_offset_in_bits = 1;
defparam ram_block3a46.data_interleave_width_in_bits = 1;
defparam ram_block3a46.init_file = "meminit.hex";
defparam ram_block3a46.init_file_layout = "port_a";
defparam ram_block3a46.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a46.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a46.operation_mode = "bidir_dual_port";
defparam ram_block3a46.port_a_address_clear = "none";
defparam ram_block3a46.port_a_address_width = 13;
defparam ram_block3a46.port_a_byte_enable_clock = "none";
defparam ram_block3a46.port_a_data_out_clear = "none";
defparam ram_block3a46.port_a_data_out_clock = "none";
defparam ram_block3a46.port_a_data_width = 1;
defparam ram_block3a46.port_a_first_address = 0;
defparam ram_block3a46.port_a_first_bit_number = 14;
defparam ram_block3a46.port_a_last_address = 8191;
defparam ram_block3a46.port_a_logical_ram_depth = 16384;
defparam ram_block3a46.port_a_logical_ram_width = 32;
defparam ram_block3a46.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_address_clear = "none";
defparam ram_block3a46.port_b_address_clock = "clock1";
defparam ram_block3a46.port_b_address_width = 13;
defparam ram_block3a46.port_b_data_in_clock = "clock1";
defparam ram_block3a46.port_b_data_out_clear = "none";
defparam ram_block3a46.port_b_data_out_clock = "none";
defparam ram_block3a46.port_b_data_width = 1;
defparam ram_block3a46.port_b_first_address = 0;
defparam ram_block3a46.port_b_first_bit_number = 14;
defparam ram_block3a46.port_b_last_address = 8191;
defparam ram_block3a46.port_b_logical_ram_depth = 16384;
defparam ram_block3a46.port_b_logical_ram_width = 32;
defparam ram_block3a46.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a46.port_b_read_enable_clock = "clock1";
defparam ram_block3a46.port_b_write_enable_clock = "clock1";
defparam ram_block3a46.ram_block_type = "M9K";
defparam ram_block3a46.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a46.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y29_N0
cycloneive_ram_block ram_block3a14(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[14]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[14]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a14_PORTADATAOUT_bus),
	.portbdataout(ram_block3a14_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a14.clk0_core_clock_enable = "ena0";
defparam ram_block3a14.clk1_core_clock_enable = "ena1";
defparam ram_block3a14.data_interleave_offset_in_bits = 1;
defparam ram_block3a14.data_interleave_width_in_bits = 1;
defparam ram_block3a14.init_file = "meminit.hex";
defparam ram_block3a14.init_file_layout = "port_a";
defparam ram_block3a14.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a14.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a14.operation_mode = "bidir_dual_port";
defparam ram_block3a14.port_a_address_clear = "none";
defparam ram_block3a14.port_a_address_width = 13;
defparam ram_block3a14.port_a_byte_enable_clock = "none";
defparam ram_block3a14.port_a_data_out_clear = "none";
defparam ram_block3a14.port_a_data_out_clock = "none";
defparam ram_block3a14.port_a_data_width = 1;
defparam ram_block3a14.port_a_first_address = 0;
defparam ram_block3a14.port_a_first_bit_number = 14;
defparam ram_block3a14.port_a_last_address = 8191;
defparam ram_block3a14.port_a_logical_ram_depth = 16384;
defparam ram_block3a14.port_a_logical_ram_width = 32;
defparam ram_block3a14.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_address_clear = "none";
defparam ram_block3a14.port_b_address_clock = "clock1";
defparam ram_block3a14.port_b_address_width = 13;
defparam ram_block3a14.port_b_data_in_clock = "clock1";
defparam ram_block3a14.port_b_data_out_clear = "none";
defparam ram_block3a14.port_b_data_out_clock = "none";
defparam ram_block3a14.port_b_data_width = 1;
defparam ram_block3a14.port_b_first_address = 0;
defparam ram_block3a14.port_b_first_bit_number = 14;
defparam ram_block3a14.port_b_last_address = 8191;
defparam ram_block3a14.port_b_logical_ram_depth = 16384;
defparam ram_block3a14.port_b_logical_ram_width = 32;
defparam ram_block3a14.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a14.port_b_read_enable_clock = "clock1";
defparam ram_block3a14.port_b_write_enable_clock = "clock1";
defparam ram_block3a14.ram_block_type = "M9K";
defparam ram_block3a14.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a14.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000204210000224A200503;
// synopsys translate_on

// Location: M9K_X37_Y29_N0
cycloneive_ram_block ram_block3a47(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a47_PORTADATAOUT_bus),
	.portbdataout(ram_block3a47_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a47.clk0_core_clock_enable = "ena0";
defparam ram_block3a47.clk1_core_clock_enable = "ena1";
defparam ram_block3a47.data_interleave_offset_in_bits = 1;
defparam ram_block3a47.data_interleave_width_in_bits = 1;
defparam ram_block3a47.init_file = "meminit.hex";
defparam ram_block3a47.init_file_layout = "port_a";
defparam ram_block3a47.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a47.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a47.operation_mode = "bidir_dual_port";
defparam ram_block3a47.port_a_address_clear = "none";
defparam ram_block3a47.port_a_address_width = 13;
defparam ram_block3a47.port_a_byte_enable_clock = "none";
defparam ram_block3a47.port_a_data_out_clear = "none";
defparam ram_block3a47.port_a_data_out_clock = "none";
defparam ram_block3a47.port_a_data_width = 1;
defparam ram_block3a47.port_a_first_address = 0;
defparam ram_block3a47.port_a_first_bit_number = 15;
defparam ram_block3a47.port_a_last_address = 8191;
defparam ram_block3a47.port_a_logical_ram_depth = 16384;
defparam ram_block3a47.port_a_logical_ram_width = 32;
defparam ram_block3a47.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_address_clear = "none";
defparam ram_block3a47.port_b_address_clock = "clock1";
defparam ram_block3a47.port_b_address_width = 13;
defparam ram_block3a47.port_b_data_in_clock = "clock1";
defparam ram_block3a47.port_b_data_out_clear = "none";
defparam ram_block3a47.port_b_data_out_clock = "none";
defparam ram_block3a47.port_b_data_width = 1;
defparam ram_block3a47.port_b_first_address = 0;
defparam ram_block3a47.port_b_first_bit_number = 15;
defparam ram_block3a47.port_b_last_address = 8191;
defparam ram_block3a47.port_b_logical_ram_depth = 16384;
defparam ram_block3a47.port_b_logical_ram_width = 32;
defparam ram_block3a47.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a47.port_b_read_enable_clock = "clock1";
defparam ram_block3a47.port_b_write_enable_clock = "clock1";
defparam ram_block3a47.ram_block_type = "M9K";
defparam ram_block3a47.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a47.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y35_N0
cycloneive_ram_block ram_block3a15(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[15]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[15]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a15_PORTADATAOUT_bus),
	.portbdataout(ram_block3a15_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a15.clk0_core_clock_enable = "ena0";
defparam ram_block3a15.clk1_core_clock_enable = "ena1";
defparam ram_block3a15.data_interleave_offset_in_bits = 1;
defparam ram_block3a15.data_interleave_width_in_bits = 1;
defparam ram_block3a15.init_file = "meminit.hex";
defparam ram_block3a15.init_file_layout = "port_a";
defparam ram_block3a15.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a15.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a15.operation_mode = "bidir_dual_port";
defparam ram_block3a15.port_a_address_clear = "none";
defparam ram_block3a15.port_a_address_width = 13;
defparam ram_block3a15.port_a_byte_enable_clock = "none";
defparam ram_block3a15.port_a_data_out_clear = "none";
defparam ram_block3a15.port_a_data_out_clock = "none";
defparam ram_block3a15.port_a_data_width = 1;
defparam ram_block3a15.port_a_first_address = 0;
defparam ram_block3a15.port_a_first_bit_number = 15;
defparam ram_block3a15.port_a_last_address = 8191;
defparam ram_block3a15.port_a_logical_ram_depth = 16384;
defparam ram_block3a15.port_a_logical_ram_width = 32;
defparam ram_block3a15.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_address_clear = "none";
defparam ram_block3a15.port_b_address_clock = "clock1";
defparam ram_block3a15.port_b_address_width = 13;
defparam ram_block3a15.port_b_data_in_clock = "clock1";
defparam ram_block3a15.port_b_data_out_clear = "none";
defparam ram_block3a15.port_b_data_out_clock = "none";
defparam ram_block3a15.port_b_data_width = 1;
defparam ram_block3a15.port_b_first_address = 0;
defparam ram_block3a15.port_b_first_bit_number = 15;
defparam ram_block3a15.port_b_last_address = 8191;
defparam ram_block3a15.port_b_logical_ram_depth = 16384;
defparam ram_block3a15.port_b_logical_ram_width = 32;
defparam ram_block3a15.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a15.port_b_read_enable_clock = "clock1";
defparam ram_block3a15.port_b_write_enable_clock = "clock1";
defparam ram_block3a15.ram_block_type = "M9K";
defparam ram_block3a15.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a15.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002042100002242206063;
// synopsys translate_on

// Location: M9K_X51_Y37_N0
cycloneive_ram_block ram_block3a48(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a48_PORTADATAOUT_bus),
	.portbdataout(ram_block3a48_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a48.clk0_core_clock_enable = "ena0";
defparam ram_block3a48.clk1_core_clock_enable = "ena1";
defparam ram_block3a48.data_interleave_offset_in_bits = 1;
defparam ram_block3a48.data_interleave_width_in_bits = 1;
defparam ram_block3a48.init_file = "meminit.hex";
defparam ram_block3a48.init_file_layout = "port_a";
defparam ram_block3a48.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a48.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a48.operation_mode = "bidir_dual_port";
defparam ram_block3a48.port_a_address_clear = "none";
defparam ram_block3a48.port_a_address_width = 13;
defparam ram_block3a48.port_a_byte_enable_clock = "none";
defparam ram_block3a48.port_a_data_out_clear = "none";
defparam ram_block3a48.port_a_data_out_clock = "none";
defparam ram_block3a48.port_a_data_width = 1;
defparam ram_block3a48.port_a_first_address = 0;
defparam ram_block3a48.port_a_first_bit_number = 16;
defparam ram_block3a48.port_a_last_address = 8191;
defparam ram_block3a48.port_a_logical_ram_depth = 16384;
defparam ram_block3a48.port_a_logical_ram_width = 32;
defparam ram_block3a48.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_address_clear = "none";
defparam ram_block3a48.port_b_address_clock = "clock1";
defparam ram_block3a48.port_b_address_width = 13;
defparam ram_block3a48.port_b_data_in_clock = "clock1";
defparam ram_block3a48.port_b_data_out_clear = "none";
defparam ram_block3a48.port_b_data_out_clock = "none";
defparam ram_block3a48.port_b_data_width = 1;
defparam ram_block3a48.port_b_first_address = 0;
defparam ram_block3a48.port_b_first_bit_number = 16;
defparam ram_block3a48.port_b_last_address = 8191;
defparam ram_block3a48.port_b_logical_ram_depth = 16384;
defparam ram_block3a48.port_b_logical_ram_width = 32;
defparam ram_block3a48.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a48.port_b_read_enable_clock = "clock1";
defparam ram_block3a48.port_b_write_enable_clock = "clock1";
defparam ram_block3a48.ram_block_type = "M9K";
defparam ram_block3a48.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a48.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y32_N0
cycloneive_ram_block ram_block3a16(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[16]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[16]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a16_PORTADATAOUT_bus),
	.portbdataout(ram_block3a16_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a16.clk0_core_clock_enable = "ena0";
defparam ram_block3a16.clk1_core_clock_enable = "ena1";
defparam ram_block3a16.data_interleave_offset_in_bits = 1;
defparam ram_block3a16.data_interleave_width_in_bits = 1;
defparam ram_block3a16.init_file = "meminit.hex";
defparam ram_block3a16.init_file_layout = "port_a";
defparam ram_block3a16.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a16.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a16.operation_mode = "bidir_dual_port";
defparam ram_block3a16.port_a_address_clear = "none";
defparam ram_block3a16.port_a_address_width = 13;
defparam ram_block3a16.port_a_byte_enable_clock = "none";
defparam ram_block3a16.port_a_data_out_clear = "none";
defparam ram_block3a16.port_a_data_out_clock = "none";
defparam ram_block3a16.port_a_data_width = 1;
defparam ram_block3a16.port_a_first_address = 0;
defparam ram_block3a16.port_a_first_bit_number = 16;
defparam ram_block3a16.port_a_last_address = 8191;
defparam ram_block3a16.port_a_logical_ram_depth = 16384;
defparam ram_block3a16.port_a_logical_ram_width = 32;
defparam ram_block3a16.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_address_clear = "none";
defparam ram_block3a16.port_b_address_clock = "clock1";
defparam ram_block3a16.port_b_address_width = 13;
defparam ram_block3a16.port_b_data_in_clock = "clock1";
defparam ram_block3a16.port_b_data_out_clear = "none";
defparam ram_block3a16.port_b_data_out_clock = "none";
defparam ram_block3a16.port_b_data_width = 1;
defparam ram_block3a16.port_b_first_address = 0;
defparam ram_block3a16.port_b_first_bit_number = 16;
defparam ram_block3a16.port_b_last_address = 8191;
defparam ram_block3a16.port_b_logical_ram_depth = 16384;
defparam ram_block3a16.port_b_logical_ram_width = 32;
defparam ram_block3a16.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a16.port_b_read_enable_clock = "clock1";
defparam ram_block3a16.port_b_write_enable_clock = "clock1";
defparam ram_block3a16.ram_block_type = "M9K";
defparam ram_block3a16.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a16.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000205A122003613254042;
// synopsys translate_on

// Location: M9K_X64_Y35_N0
cycloneive_ram_block ram_block3a49(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a49_PORTADATAOUT_bus),
	.portbdataout(ram_block3a49_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a49.clk0_core_clock_enable = "ena0";
defparam ram_block3a49.clk1_core_clock_enable = "ena1";
defparam ram_block3a49.data_interleave_offset_in_bits = 1;
defparam ram_block3a49.data_interleave_width_in_bits = 1;
defparam ram_block3a49.init_file = "meminit.hex";
defparam ram_block3a49.init_file_layout = "port_a";
defparam ram_block3a49.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a49.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a49.operation_mode = "bidir_dual_port";
defparam ram_block3a49.port_a_address_clear = "none";
defparam ram_block3a49.port_a_address_width = 13;
defparam ram_block3a49.port_a_byte_enable_clock = "none";
defparam ram_block3a49.port_a_data_out_clear = "none";
defparam ram_block3a49.port_a_data_out_clock = "none";
defparam ram_block3a49.port_a_data_width = 1;
defparam ram_block3a49.port_a_first_address = 0;
defparam ram_block3a49.port_a_first_bit_number = 17;
defparam ram_block3a49.port_a_last_address = 8191;
defparam ram_block3a49.port_a_logical_ram_depth = 16384;
defparam ram_block3a49.port_a_logical_ram_width = 32;
defparam ram_block3a49.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_address_clear = "none";
defparam ram_block3a49.port_b_address_clock = "clock1";
defparam ram_block3a49.port_b_address_width = 13;
defparam ram_block3a49.port_b_data_in_clock = "clock1";
defparam ram_block3a49.port_b_data_out_clear = "none";
defparam ram_block3a49.port_b_data_out_clock = "none";
defparam ram_block3a49.port_b_data_width = 1;
defparam ram_block3a49.port_b_first_address = 0;
defparam ram_block3a49.port_b_first_bit_number = 17;
defparam ram_block3a49.port_b_last_address = 8191;
defparam ram_block3a49.port_b_logical_ram_depth = 16384;
defparam ram_block3a49.port_b_logical_ram_width = 32;
defparam ram_block3a49.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a49.port_b_read_enable_clock = "clock1";
defparam ram_block3a49.port_b_write_enable_clock = "clock1";
defparam ram_block3a49.ram_block_type = "M9K";
defparam ram_block3a49.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a49.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y36_N0
cycloneive_ram_block ram_block3a17(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[17]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[17]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a17_PORTADATAOUT_bus),
	.portbdataout(ram_block3a17_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a17.clk0_core_clock_enable = "ena0";
defparam ram_block3a17.clk1_core_clock_enable = "ena1";
defparam ram_block3a17.data_interleave_offset_in_bits = 1;
defparam ram_block3a17.data_interleave_width_in_bits = 1;
defparam ram_block3a17.init_file = "meminit.hex";
defparam ram_block3a17.init_file_layout = "port_a";
defparam ram_block3a17.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a17.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a17.operation_mode = "bidir_dual_port";
defparam ram_block3a17.port_a_address_clear = "none";
defparam ram_block3a17.port_a_address_width = 13;
defparam ram_block3a17.port_a_byte_enable_clock = "none";
defparam ram_block3a17.port_a_data_out_clear = "none";
defparam ram_block3a17.port_a_data_out_clock = "none";
defparam ram_block3a17.port_a_data_width = 1;
defparam ram_block3a17.port_a_first_address = 0;
defparam ram_block3a17.port_a_first_bit_number = 17;
defparam ram_block3a17.port_a_last_address = 8191;
defparam ram_block3a17.port_a_logical_ram_depth = 16384;
defparam ram_block3a17.port_a_logical_ram_width = 32;
defparam ram_block3a17.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_address_clear = "none";
defparam ram_block3a17.port_b_address_clock = "clock1";
defparam ram_block3a17.port_b_address_width = 13;
defparam ram_block3a17.port_b_data_in_clock = "clock1";
defparam ram_block3a17.port_b_data_out_clear = "none";
defparam ram_block3a17.port_b_data_out_clock = "none";
defparam ram_block3a17.port_b_data_width = 1;
defparam ram_block3a17.port_b_first_address = 0;
defparam ram_block3a17.port_b_first_bit_number = 17;
defparam ram_block3a17.port_b_last_address = 8191;
defparam ram_block3a17.port_b_logical_ram_depth = 16384;
defparam ram_block3a17.port_b_logical_ram_width = 32;
defparam ram_block3a17.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a17.port_b_read_enable_clock = "clock1";
defparam ram_block3a17.port_b_write_enable_clock = "clock1";
defparam ram_block3a17.ram_block_type = "M9K";
defparam ram_block3a17.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a17.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000006C0340C001602060001;
// synopsys translate_on

// Location: M9K_X37_Y33_N0
cycloneive_ram_block ram_block3a50(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a50_PORTADATAOUT_bus),
	.portbdataout(ram_block3a50_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a50.clk0_core_clock_enable = "ena0";
defparam ram_block3a50.clk1_core_clock_enable = "ena1";
defparam ram_block3a50.data_interleave_offset_in_bits = 1;
defparam ram_block3a50.data_interleave_width_in_bits = 1;
defparam ram_block3a50.init_file = "meminit.hex";
defparam ram_block3a50.init_file_layout = "port_a";
defparam ram_block3a50.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a50.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a50.operation_mode = "bidir_dual_port";
defparam ram_block3a50.port_a_address_clear = "none";
defparam ram_block3a50.port_a_address_width = 13;
defparam ram_block3a50.port_a_byte_enable_clock = "none";
defparam ram_block3a50.port_a_data_out_clear = "none";
defparam ram_block3a50.port_a_data_out_clock = "none";
defparam ram_block3a50.port_a_data_width = 1;
defparam ram_block3a50.port_a_first_address = 0;
defparam ram_block3a50.port_a_first_bit_number = 18;
defparam ram_block3a50.port_a_last_address = 8191;
defparam ram_block3a50.port_a_logical_ram_depth = 16384;
defparam ram_block3a50.port_a_logical_ram_width = 32;
defparam ram_block3a50.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_address_clear = "none";
defparam ram_block3a50.port_b_address_clock = "clock1";
defparam ram_block3a50.port_b_address_width = 13;
defparam ram_block3a50.port_b_data_in_clock = "clock1";
defparam ram_block3a50.port_b_data_out_clear = "none";
defparam ram_block3a50.port_b_data_out_clock = "none";
defparam ram_block3a50.port_b_data_width = 1;
defparam ram_block3a50.port_b_first_address = 0;
defparam ram_block3a50.port_b_first_bit_number = 18;
defparam ram_block3a50.port_b_last_address = 8191;
defparam ram_block3a50.port_b_logical_ram_depth = 16384;
defparam ram_block3a50.port_b_logical_ram_width = 32;
defparam ram_block3a50.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a50.port_b_read_enable_clock = "clock1";
defparam ram_block3a50.port_b_write_enable_clock = "clock1";
defparam ram_block3a50.ram_block_type = "M9K";
defparam ram_block3a50.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a50.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y34_N0
cycloneive_ram_block ram_block3a18(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[18]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[18]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a18_PORTADATAOUT_bus),
	.portbdataout(ram_block3a18_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a18.clk0_core_clock_enable = "ena0";
defparam ram_block3a18.clk1_core_clock_enable = "ena1";
defparam ram_block3a18.data_interleave_offset_in_bits = 1;
defparam ram_block3a18.data_interleave_width_in_bits = 1;
defparam ram_block3a18.init_file = "meminit.hex";
defparam ram_block3a18.init_file_layout = "port_a";
defparam ram_block3a18.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a18.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a18.operation_mode = "bidir_dual_port";
defparam ram_block3a18.port_a_address_clear = "none";
defparam ram_block3a18.port_a_address_width = 13;
defparam ram_block3a18.port_a_byte_enable_clock = "none";
defparam ram_block3a18.port_a_data_out_clear = "none";
defparam ram_block3a18.port_a_data_out_clock = "none";
defparam ram_block3a18.port_a_data_width = 1;
defparam ram_block3a18.port_a_first_address = 0;
defparam ram_block3a18.port_a_first_bit_number = 18;
defparam ram_block3a18.port_a_last_address = 8191;
defparam ram_block3a18.port_a_logical_ram_depth = 16384;
defparam ram_block3a18.port_a_logical_ram_width = 32;
defparam ram_block3a18.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_address_clear = "none";
defparam ram_block3a18.port_b_address_clock = "clock1";
defparam ram_block3a18.port_b_address_width = 13;
defparam ram_block3a18.port_b_data_in_clock = "clock1";
defparam ram_block3a18.port_b_data_out_clear = "none";
defparam ram_block3a18.port_b_data_out_clock = "none";
defparam ram_block3a18.port_b_data_width = 1;
defparam ram_block3a18.port_b_first_address = 0;
defparam ram_block3a18.port_b_first_bit_number = 18;
defparam ram_block3a18.port_b_last_address = 8191;
defparam ram_block3a18.port_b_logical_ram_depth = 16384;
defparam ram_block3a18.port_b_logical_ram_width = 32;
defparam ram_block3a18.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a18.port_b_read_enable_clock = "clock1";
defparam ram_block3a18.port_b_write_enable_clock = "clock1";
defparam ram_block3a18.ram_block_type = "M9K";
defparam ram_block3a18.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a18.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000060C3180001703286867;
// synopsys translate_on

// Location: M9K_X64_Y31_N0
cycloneive_ram_block ram_block3a51(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a51_PORTADATAOUT_bus),
	.portbdataout(ram_block3a51_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a51.clk0_core_clock_enable = "ena0";
defparam ram_block3a51.clk1_core_clock_enable = "ena1";
defparam ram_block3a51.data_interleave_offset_in_bits = 1;
defparam ram_block3a51.data_interleave_width_in_bits = 1;
defparam ram_block3a51.init_file = "meminit.hex";
defparam ram_block3a51.init_file_layout = "port_a";
defparam ram_block3a51.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a51.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a51.operation_mode = "bidir_dual_port";
defparam ram_block3a51.port_a_address_clear = "none";
defparam ram_block3a51.port_a_address_width = 13;
defparam ram_block3a51.port_a_byte_enable_clock = "none";
defparam ram_block3a51.port_a_data_out_clear = "none";
defparam ram_block3a51.port_a_data_out_clock = "none";
defparam ram_block3a51.port_a_data_width = 1;
defparam ram_block3a51.port_a_first_address = 0;
defparam ram_block3a51.port_a_first_bit_number = 19;
defparam ram_block3a51.port_a_last_address = 8191;
defparam ram_block3a51.port_a_logical_ram_depth = 16384;
defparam ram_block3a51.port_a_logical_ram_width = 32;
defparam ram_block3a51.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_address_clear = "none";
defparam ram_block3a51.port_b_address_clock = "clock1";
defparam ram_block3a51.port_b_address_width = 13;
defparam ram_block3a51.port_b_data_in_clock = "clock1";
defparam ram_block3a51.port_b_data_out_clear = "none";
defparam ram_block3a51.port_b_data_out_clock = "none";
defparam ram_block3a51.port_b_data_width = 1;
defparam ram_block3a51.port_b_first_address = 0;
defparam ram_block3a51.port_b_first_bit_number = 19;
defparam ram_block3a51.port_b_last_address = 8191;
defparam ram_block3a51.port_b_logical_ram_depth = 16384;
defparam ram_block3a51.port_b_logical_ram_width = 32;
defparam ram_block3a51.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a51.port_b_read_enable_clock = "clock1";
defparam ram_block3a51.port_b_write_enable_clock = "clock1";
defparam ram_block3a51.ram_block_type = "M9K";
defparam ram_block3a51.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a51.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y30_N0
cycloneive_ram_block ram_block3a19(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[19]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[19]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a19_PORTADATAOUT_bus),
	.portbdataout(ram_block3a19_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a19.clk0_core_clock_enable = "ena0";
defparam ram_block3a19.clk1_core_clock_enable = "ena1";
defparam ram_block3a19.data_interleave_offset_in_bits = 1;
defparam ram_block3a19.data_interleave_width_in_bits = 1;
defparam ram_block3a19.init_file = "meminit.hex";
defparam ram_block3a19.init_file_layout = "port_a";
defparam ram_block3a19.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a19.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a19.operation_mode = "bidir_dual_port";
defparam ram_block3a19.port_a_address_clear = "none";
defparam ram_block3a19.port_a_address_width = 13;
defparam ram_block3a19.port_a_byte_enable_clock = "none";
defparam ram_block3a19.port_a_data_out_clear = "none";
defparam ram_block3a19.port_a_data_out_clock = "none";
defparam ram_block3a19.port_a_data_width = 1;
defparam ram_block3a19.port_a_first_address = 0;
defparam ram_block3a19.port_a_first_bit_number = 19;
defparam ram_block3a19.port_a_last_address = 8191;
defparam ram_block3a19.port_a_logical_ram_depth = 16384;
defparam ram_block3a19.port_a_logical_ram_width = 32;
defparam ram_block3a19.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_address_clear = "none";
defparam ram_block3a19.port_b_address_clock = "clock1";
defparam ram_block3a19.port_b_address_width = 13;
defparam ram_block3a19.port_b_data_in_clock = "clock1";
defparam ram_block3a19.port_b_data_out_clear = "none";
defparam ram_block3a19.port_b_data_out_clock = "none";
defparam ram_block3a19.port_b_data_width = 1;
defparam ram_block3a19.port_b_first_address = 0;
defparam ram_block3a19.port_b_first_bit_number = 19;
defparam ram_block3a19.port_b_last_address = 8191;
defparam ram_block3a19.port_b_logical_ram_depth = 16384;
defparam ram_block3a19.port_b_logical_ram_width = 32;
defparam ram_block3a19.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a19.port_b_read_enable_clock = "clock1";
defparam ram_block3a19.port_b_write_enable_clock = "clock1";
defparam ram_block3a19.ram_block_type = "M9K";
defparam ram_block3a19.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a19.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001C38C6E09B6D7701203;
// synopsys translate_on

// Location: M9K_X51_Y34_N0
cycloneive_ram_block ram_block3a52(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a52_PORTADATAOUT_bus),
	.portbdataout(ram_block3a52_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a52.clk0_core_clock_enable = "ena0";
defparam ram_block3a52.clk1_core_clock_enable = "ena1";
defparam ram_block3a52.data_interleave_offset_in_bits = 1;
defparam ram_block3a52.data_interleave_width_in_bits = 1;
defparam ram_block3a52.init_file = "meminit.hex";
defparam ram_block3a52.init_file_layout = "port_a";
defparam ram_block3a52.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a52.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a52.operation_mode = "bidir_dual_port";
defparam ram_block3a52.port_a_address_clear = "none";
defparam ram_block3a52.port_a_address_width = 13;
defparam ram_block3a52.port_a_byte_enable_clock = "none";
defparam ram_block3a52.port_a_data_out_clear = "none";
defparam ram_block3a52.port_a_data_out_clock = "none";
defparam ram_block3a52.port_a_data_width = 1;
defparam ram_block3a52.port_a_first_address = 0;
defparam ram_block3a52.port_a_first_bit_number = 20;
defparam ram_block3a52.port_a_last_address = 8191;
defparam ram_block3a52.port_a_logical_ram_depth = 16384;
defparam ram_block3a52.port_a_logical_ram_width = 32;
defparam ram_block3a52.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_address_clear = "none";
defparam ram_block3a52.port_b_address_clock = "clock1";
defparam ram_block3a52.port_b_address_width = 13;
defparam ram_block3a52.port_b_data_in_clock = "clock1";
defparam ram_block3a52.port_b_data_out_clear = "none";
defparam ram_block3a52.port_b_data_out_clock = "none";
defparam ram_block3a52.port_b_data_width = 1;
defparam ram_block3a52.port_b_first_address = 0;
defparam ram_block3a52.port_b_first_bit_number = 20;
defparam ram_block3a52.port_b_last_address = 8191;
defparam ram_block3a52.port_b_logical_ram_depth = 16384;
defparam ram_block3a52.port_b_logical_ram_width = 32;
defparam ram_block3a52.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a52.port_b_read_enable_clock = "clock1";
defparam ram_block3a52.port_b_write_enable_clock = "clock1";
defparam ram_block3a52.ram_block_type = "M9K";
defparam ram_block3a52.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a52.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y33_N0
cycloneive_ram_block ram_block3a20(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[20]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[20]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a20_PORTADATAOUT_bus),
	.portbdataout(ram_block3a20_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a20.clk0_core_clock_enable = "ena0";
defparam ram_block3a20.clk1_core_clock_enable = "ena1";
defparam ram_block3a20.data_interleave_offset_in_bits = 1;
defparam ram_block3a20.data_interleave_width_in_bits = 1;
defparam ram_block3a20.init_file = "meminit.hex";
defparam ram_block3a20.init_file_layout = "port_a";
defparam ram_block3a20.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a20.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a20.operation_mode = "bidir_dual_port";
defparam ram_block3a20.port_a_address_clear = "none";
defparam ram_block3a20.port_a_address_width = 13;
defparam ram_block3a20.port_a_byte_enable_clock = "none";
defparam ram_block3a20.port_a_data_out_clear = "none";
defparam ram_block3a20.port_a_data_out_clock = "none";
defparam ram_block3a20.port_a_data_width = 1;
defparam ram_block3a20.port_a_first_address = 0;
defparam ram_block3a20.port_a_first_bit_number = 20;
defparam ram_block3a20.port_a_last_address = 8191;
defparam ram_block3a20.port_a_logical_ram_depth = 16384;
defparam ram_block3a20.port_a_logical_ram_width = 32;
defparam ram_block3a20.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_address_clear = "none";
defparam ram_block3a20.port_b_address_clock = "clock1";
defparam ram_block3a20.port_b_address_width = 13;
defparam ram_block3a20.port_b_data_in_clock = "clock1";
defparam ram_block3a20.port_b_data_out_clear = "none";
defparam ram_block3a20.port_b_data_out_clock = "none";
defparam ram_block3a20.port_b_data_width = 1;
defparam ram_block3a20.port_b_first_address = 0;
defparam ram_block3a20.port_b_first_bit_number = 20;
defparam ram_block3a20.port_b_last_address = 8191;
defparam ram_block3a20.port_b_logical_ram_depth = 16384;
defparam ram_block3a20.port_b_logical_ram_width = 32;
defparam ram_block3a20.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a20.port_b_read_enable_clock = "clock1";
defparam ram_block3a20.port_b_write_enable_clock = "clock1";
defparam ram_block3a20.ram_block_type = "M9K";
defparam ram_block3a20.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a20.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000A0832F000B;
// synopsys translate_on

// Location: M9K_X64_Y37_N0
cycloneive_ram_block ram_block3a53(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a53_PORTADATAOUT_bus),
	.portbdataout(ram_block3a53_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a53.clk0_core_clock_enable = "ena0";
defparam ram_block3a53.clk1_core_clock_enable = "ena1";
defparam ram_block3a53.data_interleave_offset_in_bits = 1;
defparam ram_block3a53.data_interleave_width_in_bits = 1;
defparam ram_block3a53.init_file = "meminit.hex";
defparam ram_block3a53.init_file_layout = "port_a";
defparam ram_block3a53.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a53.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a53.operation_mode = "bidir_dual_port";
defparam ram_block3a53.port_a_address_clear = "none";
defparam ram_block3a53.port_a_address_width = 13;
defparam ram_block3a53.port_a_byte_enable_clock = "none";
defparam ram_block3a53.port_a_data_out_clear = "none";
defparam ram_block3a53.port_a_data_out_clock = "none";
defparam ram_block3a53.port_a_data_width = 1;
defparam ram_block3a53.port_a_first_address = 0;
defparam ram_block3a53.port_a_first_bit_number = 21;
defparam ram_block3a53.port_a_last_address = 8191;
defparam ram_block3a53.port_a_logical_ram_depth = 16384;
defparam ram_block3a53.port_a_logical_ram_width = 32;
defparam ram_block3a53.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_address_clear = "none";
defparam ram_block3a53.port_b_address_clock = "clock1";
defparam ram_block3a53.port_b_address_width = 13;
defparam ram_block3a53.port_b_data_in_clock = "clock1";
defparam ram_block3a53.port_b_data_out_clear = "none";
defparam ram_block3a53.port_b_data_out_clock = "none";
defparam ram_block3a53.port_b_data_width = 1;
defparam ram_block3a53.port_b_first_address = 0;
defparam ram_block3a53.port_b_first_bit_number = 21;
defparam ram_block3a53.port_b_last_address = 8191;
defparam ram_block3a53.port_b_logical_ram_depth = 16384;
defparam ram_block3a53.port_b_logical_ram_width = 32;
defparam ram_block3a53.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a53.port_b_read_enable_clock = "clock1";
defparam ram_block3a53.port_b_write_enable_clock = "clock1";
defparam ram_block3a53.ram_block_type = "M9K";
defparam ram_block3a53.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a53.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y34_N0
cycloneive_ram_block ram_block3a21(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[21]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[21]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a21_PORTADATAOUT_bus),
	.portbdataout(ram_block3a21_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a21.clk0_core_clock_enable = "ena0";
defparam ram_block3a21.clk1_core_clock_enable = "ena1";
defparam ram_block3a21.data_interleave_offset_in_bits = 1;
defparam ram_block3a21.data_interleave_width_in_bits = 1;
defparam ram_block3a21.init_file = "meminit.hex";
defparam ram_block3a21.init_file_layout = "port_a";
defparam ram_block3a21.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a21.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a21.operation_mode = "bidir_dual_port";
defparam ram_block3a21.port_a_address_clear = "none";
defparam ram_block3a21.port_a_address_width = 13;
defparam ram_block3a21.port_a_byte_enable_clock = "none";
defparam ram_block3a21.port_a_data_out_clear = "none";
defparam ram_block3a21.port_a_data_out_clock = "none";
defparam ram_block3a21.port_a_data_width = 1;
defparam ram_block3a21.port_a_first_address = 0;
defparam ram_block3a21.port_a_first_bit_number = 21;
defparam ram_block3a21.port_a_last_address = 8191;
defparam ram_block3a21.port_a_logical_ram_depth = 16384;
defparam ram_block3a21.port_a_logical_ram_width = 32;
defparam ram_block3a21.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_address_clear = "none";
defparam ram_block3a21.port_b_address_clock = "clock1";
defparam ram_block3a21.port_b_address_width = 13;
defparam ram_block3a21.port_b_data_in_clock = "clock1";
defparam ram_block3a21.port_b_data_out_clear = "none";
defparam ram_block3a21.port_b_data_out_clock = "none";
defparam ram_block3a21.port_b_data_width = 1;
defparam ram_block3a21.port_b_first_address = 0;
defparam ram_block3a21.port_b_first_bit_number = 21;
defparam ram_block3a21.port_b_last_address = 8191;
defparam ram_block3a21.port_b_logical_ram_depth = 16384;
defparam ram_block3a21.port_b_logical_ram_width = 32;
defparam ram_block3a21.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a21.port_b_read_enable_clock = "clock1";
defparam ram_block3a21.port_b_write_enable_clock = "clock1";
defparam ram_block3a21.ram_block_type = "M9K";
defparam ram_block3a21.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a21.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002A142119BCBBAB600000;
// synopsys translate_on

// Location: M9K_X78_Y37_N0
cycloneive_ram_block ram_block3a54(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a54_PORTADATAOUT_bus),
	.portbdataout(ram_block3a54_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a54.clk0_core_clock_enable = "ena0";
defparam ram_block3a54.clk1_core_clock_enable = "ena1";
defparam ram_block3a54.data_interleave_offset_in_bits = 1;
defparam ram_block3a54.data_interleave_width_in_bits = 1;
defparam ram_block3a54.init_file = "meminit.hex";
defparam ram_block3a54.init_file_layout = "port_a";
defparam ram_block3a54.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a54.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a54.operation_mode = "bidir_dual_port";
defparam ram_block3a54.port_a_address_clear = "none";
defparam ram_block3a54.port_a_address_width = 13;
defparam ram_block3a54.port_a_byte_enable_clock = "none";
defparam ram_block3a54.port_a_data_out_clear = "none";
defparam ram_block3a54.port_a_data_out_clock = "none";
defparam ram_block3a54.port_a_data_width = 1;
defparam ram_block3a54.port_a_first_address = 0;
defparam ram_block3a54.port_a_first_bit_number = 22;
defparam ram_block3a54.port_a_last_address = 8191;
defparam ram_block3a54.port_a_logical_ram_depth = 16384;
defparam ram_block3a54.port_a_logical_ram_width = 32;
defparam ram_block3a54.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_address_clear = "none";
defparam ram_block3a54.port_b_address_clock = "clock1";
defparam ram_block3a54.port_b_address_width = 13;
defparam ram_block3a54.port_b_data_in_clock = "clock1";
defparam ram_block3a54.port_b_data_out_clear = "none";
defparam ram_block3a54.port_b_data_out_clock = "none";
defparam ram_block3a54.port_b_data_width = 1;
defparam ram_block3a54.port_b_first_address = 0;
defparam ram_block3a54.port_b_first_bit_number = 22;
defparam ram_block3a54.port_b_last_address = 8191;
defparam ram_block3a54.port_b_logical_ram_depth = 16384;
defparam ram_block3a54.port_b_logical_ram_width = 32;
defparam ram_block3a54.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a54.port_b_read_enable_clock = "clock1";
defparam ram_block3a54.port_b_write_enable_clock = "clock1";
defparam ram_block3a54.ram_block_type = "M9K";
defparam ram_block3a54.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a54.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y36_N0
cycloneive_ram_block ram_block3a22(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[22]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[22]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a22_PORTADATAOUT_bus),
	.portbdataout(ram_block3a22_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a22.clk0_core_clock_enable = "ena0";
defparam ram_block3a22.clk1_core_clock_enable = "ena1";
defparam ram_block3a22.data_interleave_offset_in_bits = 1;
defparam ram_block3a22.data_interleave_width_in_bits = 1;
defparam ram_block3a22.init_file = "meminit.hex";
defparam ram_block3a22.init_file_layout = "port_a";
defparam ram_block3a22.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a22.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a22.operation_mode = "bidir_dual_port";
defparam ram_block3a22.port_a_address_clear = "none";
defparam ram_block3a22.port_a_address_width = 13;
defparam ram_block3a22.port_a_byte_enable_clock = "none";
defparam ram_block3a22.port_a_data_out_clear = "none";
defparam ram_block3a22.port_a_data_out_clock = "none";
defparam ram_block3a22.port_a_data_width = 1;
defparam ram_block3a22.port_a_first_address = 0;
defparam ram_block3a22.port_a_first_bit_number = 22;
defparam ram_block3a22.port_a_last_address = 8191;
defparam ram_block3a22.port_a_logical_ram_depth = 16384;
defparam ram_block3a22.port_a_logical_ram_width = 32;
defparam ram_block3a22.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_address_clear = "none";
defparam ram_block3a22.port_b_address_clock = "clock1";
defparam ram_block3a22.port_b_address_width = 13;
defparam ram_block3a22.port_b_data_in_clock = "clock1";
defparam ram_block3a22.port_b_data_out_clear = "none";
defparam ram_block3a22.port_b_data_out_clock = "none";
defparam ram_block3a22.port_b_data_width = 1;
defparam ram_block3a22.port_b_first_address = 0;
defparam ram_block3a22.port_b_first_bit_number = 22;
defparam ram_block3a22.port_b_last_address = 8191;
defparam ram_block3a22.port_b_logical_ram_depth = 16384;
defparam ram_block3a22.port_b_logical_ram_width = 32;
defparam ram_block3a22.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a22.port_b_read_enable_clock = "clock1";
defparam ram_block3a22.port_b_write_enable_clock = "clock1";
defparam ram_block3a22.ram_block_type = "M9K";
defparam ram_block3a22.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a22.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E403004A40002000000;
// synopsys translate_on

// Location: M9K_X64_Y33_N0
cycloneive_ram_block ram_block3a55(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a55_PORTADATAOUT_bus),
	.portbdataout(ram_block3a55_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a55.clk0_core_clock_enable = "ena0";
defparam ram_block3a55.clk1_core_clock_enable = "ena1";
defparam ram_block3a55.data_interleave_offset_in_bits = 1;
defparam ram_block3a55.data_interleave_width_in_bits = 1;
defparam ram_block3a55.init_file = "meminit.hex";
defparam ram_block3a55.init_file_layout = "port_a";
defparam ram_block3a55.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a55.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a55.operation_mode = "bidir_dual_port";
defparam ram_block3a55.port_a_address_clear = "none";
defparam ram_block3a55.port_a_address_width = 13;
defparam ram_block3a55.port_a_byte_enable_clock = "none";
defparam ram_block3a55.port_a_data_out_clear = "none";
defparam ram_block3a55.port_a_data_out_clock = "none";
defparam ram_block3a55.port_a_data_width = 1;
defparam ram_block3a55.port_a_first_address = 0;
defparam ram_block3a55.port_a_first_bit_number = 23;
defparam ram_block3a55.port_a_last_address = 8191;
defparam ram_block3a55.port_a_logical_ram_depth = 16384;
defparam ram_block3a55.port_a_logical_ram_width = 32;
defparam ram_block3a55.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_address_clear = "none";
defparam ram_block3a55.port_b_address_clock = "clock1";
defparam ram_block3a55.port_b_address_width = 13;
defparam ram_block3a55.port_b_data_in_clock = "clock1";
defparam ram_block3a55.port_b_data_out_clear = "none";
defparam ram_block3a55.port_b_data_out_clock = "none";
defparam ram_block3a55.port_b_data_width = 1;
defparam ram_block3a55.port_b_first_address = 0;
defparam ram_block3a55.port_b_first_bit_number = 23;
defparam ram_block3a55.port_b_last_address = 8191;
defparam ram_block3a55.port_b_logical_ram_depth = 16384;
defparam ram_block3a55.port_b_logical_ram_width = 32;
defparam ram_block3a55.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a55.port_b_read_enable_clock = "clock1";
defparam ram_block3a55.port_b_write_enable_clock = "clock1";
defparam ram_block3a55.ram_block_type = "M9K";
defparam ram_block3a55.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a55.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y32_N0
cycloneive_ram_block ram_block3a23(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[23]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[23]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a23_PORTADATAOUT_bus),
	.portbdataout(ram_block3a23_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a23.clk0_core_clock_enable = "ena0";
defparam ram_block3a23.clk1_core_clock_enable = "ena1";
defparam ram_block3a23.data_interleave_offset_in_bits = 1;
defparam ram_block3a23.data_interleave_width_in_bits = 1;
defparam ram_block3a23.init_file = "meminit.hex";
defparam ram_block3a23.init_file_layout = "port_a";
defparam ram_block3a23.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a23.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a23.operation_mode = "bidir_dual_port";
defparam ram_block3a23.port_a_address_clear = "none";
defparam ram_block3a23.port_a_address_width = 13;
defparam ram_block3a23.port_a_byte_enable_clock = "none";
defparam ram_block3a23.port_a_data_out_clear = "none";
defparam ram_block3a23.port_a_data_out_clock = "none";
defparam ram_block3a23.port_a_data_width = 1;
defparam ram_block3a23.port_a_first_address = 0;
defparam ram_block3a23.port_a_first_bit_number = 23;
defparam ram_block3a23.port_a_last_address = 8191;
defparam ram_block3a23.port_a_logical_ram_depth = 16384;
defparam ram_block3a23.port_a_logical_ram_width = 32;
defparam ram_block3a23.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_address_clear = "none";
defparam ram_block3a23.port_b_address_clock = "clock1";
defparam ram_block3a23.port_b_address_width = 13;
defparam ram_block3a23.port_b_data_in_clock = "clock1";
defparam ram_block3a23.port_b_data_out_clear = "none";
defparam ram_block3a23.port_b_data_out_clock = "none";
defparam ram_block3a23.port_b_data_width = 1;
defparam ram_block3a23.port_b_first_address = 0;
defparam ram_block3a23.port_b_first_bit_number = 23;
defparam ram_block3a23.port_b_last_address = 8191;
defparam ram_block3a23.port_b_logical_ram_depth = 16384;
defparam ram_block3a23.port_b_logical_ram_width = 32;
defparam ram_block3a23.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a23.port_b_read_enable_clock = "clock1";
defparam ram_block3a23.port_b_write_enable_clock = "clock1";
defparam ram_block3a23.ram_block_type = "M9K";
defparam ram_block3a23.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a23.mem_init0 = 2048'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002E5CB187BC004B601000;
// synopsys translate_on

// Location: M9K_X37_Y32_N0
cycloneive_ram_block ram_block3a56(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a56_PORTADATAOUT_bus),
	.portbdataout(ram_block3a56_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a56.clk0_core_clock_enable = "ena0";
defparam ram_block3a56.clk1_core_clock_enable = "ena1";
defparam ram_block3a56.data_interleave_offset_in_bits = 1;
defparam ram_block3a56.data_interleave_width_in_bits = 1;
defparam ram_block3a56.init_file = "meminit.hex";
defparam ram_block3a56.init_file_layout = "port_a";
defparam ram_block3a56.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a56.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a56.operation_mode = "bidir_dual_port";
defparam ram_block3a56.port_a_address_clear = "none";
defparam ram_block3a56.port_a_address_width = 13;
defparam ram_block3a56.port_a_byte_enable_clock = "none";
defparam ram_block3a56.port_a_data_out_clear = "none";
defparam ram_block3a56.port_a_data_out_clock = "none";
defparam ram_block3a56.port_a_data_width = 1;
defparam ram_block3a56.port_a_first_address = 0;
defparam ram_block3a56.port_a_first_bit_number = 24;
defparam ram_block3a56.port_a_last_address = 8191;
defparam ram_block3a56.port_a_logical_ram_depth = 16384;
defparam ram_block3a56.port_a_logical_ram_width = 32;
defparam ram_block3a56.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_address_clear = "none";
defparam ram_block3a56.port_b_address_clock = "clock1";
defparam ram_block3a56.port_b_address_width = 13;
defparam ram_block3a56.port_b_data_in_clock = "clock1";
defparam ram_block3a56.port_b_data_out_clear = "none";
defparam ram_block3a56.port_b_data_out_clock = "none";
defparam ram_block3a56.port_b_data_width = 1;
defparam ram_block3a56.port_b_first_address = 0;
defparam ram_block3a56.port_b_first_bit_number = 24;
defparam ram_block3a56.port_b_last_address = 8191;
defparam ram_block3a56.port_b_logical_ram_depth = 16384;
defparam ram_block3a56.port_b_logical_ram_width = 32;
defparam ram_block3a56.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a56.port_b_read_enable_clock = "clock1";
defparam ram_block3a56.port_b_write_enable_clock = "clock1";
defparam ram_block3a56.ram_block_type = "M9K";
defparam ram_block3a56.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a56.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y36_N0
cycloneive_ram_block ram_block3a24(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[24]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[24]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a24_PORTADATAOUT_bus),
	.portbdataout(ram_block3a24_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a24.clk0_core_clock_enable = "ena0";
defparam ram_block3a24.clk1_core_clock_enable = "ena1";
defparam ram_block3a24.data_interleave_offset_in_bits = 1;
defparam ram_block3a24.data_interleave_width_in_bits = 1;
defparam ram_block3a24.init_file = "meminit.hex";
defparam ram_block3a24.init_file_layout = "port_a";
defparam ram_block3a24.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a24.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a24.operation_mode = "bidir_dual_port";
defparam ram_block3a24.port_a_address_clear = "none";
defparam ram_block3a24.port_a_address_width = 13;
defparam ram_block3a24.port_a_byte_enable_clock = "none";
defparam ram_block3a24.port_a_data_out_clear = "none";
defparam ram_block3a24.port_a_data_out_clock = "none";
defparam ram_block3a24.port_a_data_width = 1;
defparam ram_block3a24.port_a_first_address = 0;
defparam ram_block3a24.port_a_first_bit_number = 24;
defparam ram_block3a24.port_a_last_address = 8191;
defparam ram_block3a24.port_a_logical_ram_depth = 16384;
defparam ram_block3a24.port_a_logical_ram_width = 32;
defparam ram_block3a24.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_address_clear = "none";
defparam ram_block3a24.port_b_address_clock = "clock1";
defparam ram_block3a24.port_b_address_width = 13;
defparam ram_block3a24.port_b_data_in_clock = "clock1";
defparam ram_block3a24.port_b_data_out_clear = "none";
defparam ram_block3a24.port_b_data_out_clock = "none";
defparam ram_block3a24.port_b_data_width = 1;
defparam ram_block3a24.port_b_first_address = 0;
defparam ram_block3a24.port_b_first_bit_number = 24;
defparam ram_block3a24.port_b_last_address = 8191;
defparam ram_block3a24.port_b_logical_ram_depth = 16384;
defparam ram_block3a24.port_b_logical_ram_width = 32;
defparam ram_block3a24.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a24.port_b_read_enable_clock = "clock1";
defparam ram_block3a24.port_b_write_enable_clock = "clock1";
defparam ram_block3a24.ram_block_type = "M9K";
defparam ram_block3a24.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a24.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000021830C680DB793600400;
// synopsys translate_on

// Location: M9K_X51_Y30_N0
cycloneive_ram_block ram_block3a57(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a57_PORTADATAOUT_bus),
	.portbdataout(ram_block3a57_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a57.clk0_core_clock_enable = "ena0";
defparam ram_block3a57.clk1_core_clock_enable = "ena1";
defparam ram_block3a57.data_interleave_offset_in_bits = 1;
defparam ram_block3a57.data_interleave_width_in_bits = 1;
defparam ram_block3a57.init_file = "meminit.hex";
defparam ram_block3a57.init_file_layout = "port_a";
defparam ram_block3a57.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a57.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a57.operation_mode = "bidir_dual_port";
defparam ram_block3a57.port_a_address_clear = "none";
defparam ram_block3a57.port_a_address_width = 13;
defparam ram_block3a57.port_a_byte_enable_clock = "none";
defparam ram_block3a57.port_a_data_out_clear = "none";
defparam ram_block3a57.port_a_data_out_clock = "none";
defparam ram_block3a57.port_a_data_width = 1;
defparam ram_block3a57.port_a_first_address = 0;
defparam ram_block3a57.port_a_first_bit_number = 25;
defparam ram_block3a57.port_a_last_address = 8191;
defparam ram_block3a57.port_a_logical_ram_depth = 16384;
defparam ram_block3a57.port_a_logical_ram_width = 32;
defparam ram_block3a57.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_address_clear = "none";
defparam ram_block3a57.port_b_address_clock = "clock1";
defparam ram_block3a57.port_b_address_width = 13;
defparam ram_block3a57.port_b_data_in_clock = "clock1";
defparam ram_block3a57.port_b_data_out_clear = "none";
defparam ram_block3a57.port_b_data_out_clock = "none";
defparam ram_block3a57.port_b_data_width = 1;
defparam ram_block3a57.port_b_first_address = 0;
defparam ram_block3a57.port_b_first_bit_number = 25;
defparam ram_block3a57.port_b_last_address = 8191;
defparam ram_block3a57.port_b_logical_ram_depth = 16384;
defparam ram_block3a57.port_b_logical_ram_width = 32;
defparam ram_block3a57.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a57.port_b_read_enable_clock = "clock1";
defparam ram_block3a57.port_b_write_enable_clock = "clock1";
defparam ram_block3a57.ram_block_type = "M9K";
defparam ram_block3a57.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a57.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y31_N0
cycloneive_ram_block ram_block3a25(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[25]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[25]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a25_PORTADATAOUT_bus),
	.portbdataout(ram_block3a25_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a25.clk0_core_clock_enable = "ena0";
defparam ram_block3a25.clk1_core_clock_enable = "ena1";
defparam ram_block3a25.data_interleave_offset_in_bits = 1;
defparam ram_block3a25.data_interleave_width_in_bits = 1;
defparam ram_block3a25.init_file = "meminit.hex";
defparam ram_block3a25.init_file_layout = "port_a";
defparam ram_block3a25.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a25.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a25.operation_mode = "bidir_dual_port";
defparam ram_block3a25.port_a_address_clear = "none";
defparam ram_block3a25.port_a_address_width = 13;
defparam ram_block3a25.port_a_byte_enable_clock = "none";
defparam ram_block3a25.port_a_data_out_clear = "none";
defparam ram_block3a25.port_a_data_out_clock = "none";
defparam ram_block3a25.port_a_data_width = 1;
defparam ram_block3a25.port_a_first_address = 0;
defparam ram_block3a25.port_a_first_bit_number = 25;
defparam ram_block3a25.port_a_last_address = 8191;
defparam ram_block3a25.port_a_logical_ram_depth = 16384;
defparam ram_block3a25.port_a_logical_ram_width = 32;
defparam ram_block3a25.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_address_clear = "none";
defparam ram_block3a25.port_b_address_clock = "clock1";
defparam ram_block3a25.port_b_address_width = 13;
defparam ram_block3a25.port_b_data_in_clock = "clock1";
defparam ram_block3a25.port_b_data_out_clear = "none";
defparam ram_block3a25.port_b_data_out_clock = "none";
defparam ram_block3a25.port_b_data_width = 1;
defparam ram_block3a25.port_b_first_address = 0;
defparam ram_block3a25.port_b_first_bit_number = 25;
defparam ram_block3a25.port_b_last_address = 8191;
defparam ram_block3a25.port_b_logical_ram_depth = 16384;
defparam ram_block3a25.port_b_logical_ram_width = 32;
defparam ram_block3a25.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a25.port_b_read_enable_clock = "clock1";
defparam ram_block3a25.port_b_write_enable_clock = "clock1";
defparam ram_block3a25.ram_block_type = "M9K";
defparam ram_block3a25.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a25.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000200000000CB783600310;
// synopsys translate_on

// Location: M9K_X51_Y36_N0
cycloneive_ram_block ram_block3a58(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a58_PORTADATAOUT_bus),
	.portbdataout(ram_block3a58_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a58.clk0_core_clock_enable = "ena0";
defparam ram_block3a58.clk1_core_clock_enable = "ena1";
defparam ram_block3a58.data_interleave_offset_in_bits = 1;
defparam ram_block3a58.data_interleave_width_in_bits = 1;
defparam ram_block3a58.init_file = "meminit.hex";
defparam ram_block3a58.init_file_layout = "port_a";
defparam ram_block3a58.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a58.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a58.operation_mode = "bidir_dual_port";
defparam ram_block3a58.port_a_address_clear = "none";
defparam ram_block3a58.port_a_address_width = 13;
defparam ram_block3a58.port_a_byte_enable_clock = "none";
defparam ram_block3a58.port_a_data_out_clear = "none";
defparam ram_block3a58.port_a_data_out_clock = "none";
defparam ram_block3a58.port_a_data_width = 1;
defparam ram_block3a58.port_a_first_address = 0;
defparam ram_block3a58.port_a_first_bit_number = 26;
defparam ram_block3a58.port_a_last_address = 8191;
defparam ram_block3a58.port_a_logical_ram_depth = 16384;
defparam ram_block3a58.port_a_logical_ram_width = 32;
defparam ram_block3a58.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_address_clear = "none";
defparam ram_block3a58.port_b_address_clock = "clock1";
defparam ram_block3a58.port_b_address_width = 13;
defparam ram_block3a58.port_b_data_in_clock = "clock1";
defparam ram_block3a58.port_b_data_out_clear = "none";
defparam ram_block3a58.port_b_data_out_clock = "none";
defparam ram_block3a58.port_b_data_width = 1;
defparam ram_block3a58.port_b_first_address = 0;
defparam ram_block3a58.port_b_first_bit_number = 26;
defparam ram_block3a58.port_b_last_address = 8191;
defparam ram_block3a58.port_b_logical_ram_depth = 16384;
defparam ram_block3a58.port_b_logical_ram_width = 32;
defparam ram_block3a58.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a58.port_b_read_enable_clock = "clock1";
defparam ram_block3a58.port_b_write_enable_clock = "clock1";
defparam ram_block3a58.ram_block_type = "M9K";
defparam ram_block3a58.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a58.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y35_N0
cycloneive_ram_block ram_block3a26(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[26]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[26]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a26_PORTADATAOUT_bus),
	.portbdataout(ram_block3a26_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a26.clk0_core_clock_enable = "ena0";
defparam ram_block3a26.clk1_core_clock_enable = "ena1";
defparam ram_block3a26.data_interleave_offset_in_bits = 1;
defparam ram_block3a26.data_interleave_width_in_bits = 1;
defparam ram_block3a26.init_file = "meminit.hex";
defparam ram_block3a26.init_file_layout = "port_a";
defparam ram_block3a26.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a26.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a26.operation_mode = "bidir_dual_port";
defparam ram_block3a26.port_a_address_clear = "none";
defparam ram_block3a26.port_a_address_width = 13;
defparam ram_block3a26.port_a_byte_enable_clock = "none";
defparam ram_block3a26.port_a_data_out_clear = "none";
defparam ram_block3a26.port_a_data_out_clock = "none";
defparam ram_block3a26.port_a_data_width = 1;
defparam ram_block3a26.port_a_first_address = 0;
defparam ram_block3a26.port_a_first_bit_number = 26;
defparam ram_block3a26.port_a_last_address = 8191;
defparam ram_block3a26.port_a_logical_ram_depth = 16384;
defparam ram_block3a26.port_a_logical_ram_width = 32;
defparam ram_block3a26.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_address_clear = "none";
defparam ram_block3a26.port_b_address_clock = "clock1";
defparam ram_block3a26.port_b_address_width = 13;
defparam ram_block3a26.port_b_data_in_clock = "clock1";
defparam ram_block3a26.port_b_data_out_clear = "none";
defparam ram_block3a26.port_b_data_out_clock = "none";
defparam ram_block3a26.port_b_data_width = 1;
defparam ram_block3a26.port_b_first_address = 0;
defparam ram_block3a26.port_b_first_bit_number = 26;
defparam ram_block3a26.port_b_last_address = 8191;
defparam ram_block3a26.port_b_logical_ram_depth = 16384;
defparam ram_block3a26.port_b_logical_ram_width = 32;
defparam ram_block3a26.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a26.port_b_read_enable_clock = "clock1";
defparam ram_block3a26.port_b_write_enable_clock = "clock1";
defparam ram_block3a26.ram_block_type = "M9K";
defparam ram_block3a26.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a26.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000007CFBDE639B287F0888F;
// synopsys translate_on

// Location: M9K_X64_Y24_N0
cycloneive_ram_block ram_block3a59(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a59_PORTADATAOUT_bus),
	.portbdataout(ram_block3a59_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a59.clk0_core_clock_enable = "ena0";
defparam ram_block3a59.clk1_core_clock_enable = "ena1";
defparam ram_block3a59.data_interleave_offset_in_bits = 1;
defparam ram_block3a59.data_interleave_width_in_bits = 1;
defparam ram_block3a59.init_file = "meminit.hex";
defparam ram_block3a59.init_file_layout = "port_a";
defparam ram_block3a59.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a59.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a59.operation_mode = "bidir_dual_port";
defparam ram_block3a59.port_a_address_clear = "none";
defparam ram_block3a59.port_a_address_width = 13;
defparam ram_block3a59.port_a_byte_enable_clock = "none";
defparam ram_block3a59.port_a_data_out_clear = "none";
defparam ram_block3a59.port_a_data_out_clock = "none";
defparam ram_block3a59.port_a_data_width = 1;
defparam ram_block3a59.port_a_first_address = 0;
defparam ram_block3a59.port_a_first_bit_number = 27;
defparam ram_block3a59.port_a_last_address = 8191;
defparam ram_block3a59.port_a_logical_ram_depth = 16384;
defparam ram_block3a59.port_a_logical_ram_width = 32;
defparam ram_block3a59.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_address_clear = "none";
defparam ram_block3a59.port_b_address_clock = "clock1";
defparam ram_block3a59.port_b_address_width = 13;
defparam ram_block3a59.port_b_data_in_clock = "clock1";
defparam ram_block3a59.port_b_data_out_clear = "none";
defparam ram_block3a59.port_b_data_out_clock = "none";
defparam ram_block3a59.port_b_data_width = 1;
defparam ram_block3a59.port_b_first_address = 0;
defparam ram_block3a59.port_b_first_bit_number = 27;
defparam ram_block3a59.port_b_last_address = 8191;
defparam ram_block3a59.port_b_logical_ram_depth = 16384;
defparam ram_block3a59.port_b_logical_ram_width = 32;
defparam ram_block3a59.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a59.port_b_read_enable_clock = "clock1";
defparam ram_block3a59.port_b_write_enable_clock = "clock1";
defparam ram_block3a59.ram_block_type = "M9K";
defparam ram_block3a59.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a59.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X78_Y24_N0
cycloneive_ram_block ram_block3a27(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[27]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[27]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a27_PORTADATAOUT_bus),
	.portbdataout(ram_block3a27_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a27.clk0_core_clock_enable = "ena0";
defparam ram_block3a27.clk1_core_clock_enable = "ena1";
defparam ram_block3a27.data_interleave_offset_in_bits = 1;
defparam ram_block3a27.data_interleave_width_in_bits = 1;
defparam ram_block3a27.init_file = "meminit.hex";
defparam ram_block3a27.init_file_layout = "port_a";
defparam ram_block3a27.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a27.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a27.operation_mode = "bidir_dual_port";
defparam ram_block3a27.port_a_address_clear = "none";
defparam ram_block3a27.port_a_address_width = 13;
defparam ram_block3a27.port_a_byte_enable_clock = "none";
defparam ram_block3a27.port_a_data_out_clear = "none";
defparam ram_block3a27.port_a_data_out_clock = "none";
defparam ram_block3a27.port_a_data_width = 1;
defparam ram_block3a27.port_a_first_address = 0;
defparam ram_block3a27.port_a_first_bit_number = 27;
defparam ram_block3a27.port_a_last_address = 8191;
defparam ram_block3a27.port_a_logical_ram_depth = 16384;
defparam ram_block3a27.port_a_logical_ram_width = 32;
defparam ram_block3a27.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_address_clear = "none";
defparam ram_block3a27.port_b_address_clock = "clock1";
defparam ram_block3a27.port_b_address_width = 13;
defparam ram_block3a27.port_b_data_in_clock = "clock1";
defparam ram_block3a27.port_b_data_out_clear = "none";
defparam ram_block3a27.port_b_data_out_clock = "none";
defparam ram_block3a27.port_b_data_width = 1;
defparam ram_block3a27.port_b_first_address = 0;
defparam ram_block3a27.port_b_first_bit_number = 27;
defparam ram_block3a27.port_b_last_address = 8191;
defparam ram_block3a27.port_b_logical_ram_depth = 16384;
defparam ram_block3a27.port_b_logical_ram_width = 32;
defparam ram_block3a27.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a27.port_b_read_enable_clock = "clock1";
defparam ram_block3a27.port_b_write_enable_clock = "clock1";
defparam ram_block3a27.ram_block_type = "M9K";
defparam ram_block3a27.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a27.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010E1C6264AD282C08088;
// synopsys translate_on

// Location: M9K_X51_Y27_N0
cycloneive_ram_block ram_block3a60(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a60_PORTADATAOUT_bus),
	.portbdataout(ram_block3a60_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a60.clk0_core_clock_enable = "ena0";
defparam ram_block3a60.clk1_core_clock_enable = "ena1";
defparam ram_block3a60.data_interleave_offset_in_bits = 1;
defparam ram_block3a60.data_interleave_width_in_bits = 1;
defparam ram_block3a60.init_file = "meminit.hex";
defparam ram_block3a60.init_file_layout = "port_a";
defparam ram_block3a60.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a60.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a60.operation_mode = "bidir_dual_port";
defparam ram_block3a60.port_a_address_clear = "none";
defparam ram_block3a60.port_a_address_width = 13;
defparam ram_block3a60.port_a_byte_enable_clock = "none";
defparam ram_block3a60.port_a_data_out_clear = "none";
defparam ram_block3a60.port_a_data_out_clock = "none";
defparam ram_block3a60.port_a_data_width = 1;
defparam ram_block3a60.port_a_first_address = 0;
defparam ram_block3a60.port_a_first_bit_number = 28;
defparam ram_block3a60.port_a_last_address = 8191;
defparam ram_block3a60.port_a_logical_ram_depth = 16384;
defparam ram_block3a60.port_a_logical_ram_width = 32;
defparam ram_block3a60.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_address_clear = "none";
defparam ram_block3a60.port_b_address_clock = "clock1";
defparam ram_block3a60.port_b_address_width = 13;
defparam ram_block3a60.port_b_data_in_clock = "clock1";
defparam ram_block3a60.port_b_data_out_clear = "none";
defparam ram_block3a60.port_b_data_out_clock = "none";
defparam ram_block3a60.port_b_data_width = 1;
defparam ram_block3a60.port_b_first_address = 0;
defparam ram_block3a60.port_b_first_bit_number = 28;
defparam ram_block3a60.port_b_last_address = 8191;
defparam ram_block3a60.port_b_logical_ram_depth = 16384;
defparam ram_block3a60.port_b_logical_ram_width = 32;
defparam ram_block3a60.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a60.port_b_read_enable_clock = "clock1";
defparam ram_block3a60.port_b_write_enable_clock = "clock1";
defparam ram_block3a60.ram_block_type = "M9K";
defparam ram_block3a60.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a60.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y23_N0
cycloneive_ram_block ram_block3a28(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[28]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[28]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a28_PORTADATAOUT_bus),
	.portbdataout(ram_block3a28_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a28.clk0_core_clock_enable = "ena0";
defparam ram_block3a28.clk1_core_clock_enable = "ena1";
defparam ram_block3a28.data_interleave_offset_in_bits = 1;
defparam ram_block3a28.data_interleave_width_in_bits = 1;
defparam ram_block3a28.init_file = "meminit.hex";
defparam ram_block3a28.init_file_layout = "port_a";
defparam ram_block3a28.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a28.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a28.operation_mode = "bidir_dual_port";
defparam ram_block3a28.port_a_address_clear = "none";
defparam ram_block3a28.port_a_address_width = 13;
defparam ram_block3a28.port_a_byte_enable_clock = "none";
defparam ram_block3a28.port_a_data_out_clear = "none";
defparam ram_block3a28.port_a_data_out_clock = "none";
defparam ram_block3a28.port_a_data_width = 1;
defparam ram_block3a28.port_a_first_address = 0;
defparam ram_block3a28.port_a_first_bit_number = 28;
defparam ram_block3a28.port_a_last_address = 8191;
defparam ram_block3a28.port_a_logical_ram_depth = 16384;
defparam ram_block3a28.port_a_logical_ram_width = 32;
defparam ram_block3a28.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_address_clear = "none";
defparam ram_block3a28.port_b_address_clock = "clock1";
defparam ram_block3a28.port_b_address_width = 13;
defparam ram_block3a28.port_b_data_in_clock = "clock1";
defparam ram_block3a28.port_b_data_out_clear = "none";
defparam ram_block3a28.port_b_data_out_clock = "none";
defparam ram_block3a28.port_b_data_width = 1;
defparam ram_block3a28.port_b_first_address = 0;
defparam ram_block3a28.port_b_first_bit_number = 28;
defparam ram_block3a28.port_b_last_address = 8191;
defparam ram_block3a28.port_b_logical_ram_depth = 16384;
defparam ram_block3a28.port_b_logical_ram_width = 32;
defparam ram_block3a28.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a28.port_b_read_enable_clock = "clock1";
defparam ram_block3a28.port_b_write_enable_clock = "clock1";
defparam ram_block3a28.ram_block_type = "M9K";
defparam ram_block3a28.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a28.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000008100011B00926100807;
// synopsys translate_on

// Location: M9K_X37_Y30_N0
cycloneive_ram_block ram_block3a61(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a61_PORTADATAOUT_bus),
	.portbdataout(ram_block3a61_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a61.clk0_core_clock_enable = "ena0";
defparam ram_block3a61.clk1_core_clock_enable = "ena1";
defparam ram_block3a61.data_interleave_offset_in_bits = 1;
defparam ram_block3a61.data_interleave_width_in_bits = 1;
defparam ram_block3a61.init_file = "meminit.hex";
defparam ram_block3a61.init_file_layout = "port_a";
defparam ram_block3a61.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a61.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a61.operation_mode = "bidir_dual_port";
defparam ram_block3a61.port_a_address_clear = "none";
defparam ram_block3a61.port_a_address_width = 13;
defparam ram_block3a61.port_a_byte_enable_clock = "none";
defparam ram_block3a61.port_a_data_out_clear = "none";
defparam ram_block3a61.port_a_data_out_clock = "none";
defparam ram_block3a61.port_a_data_width = 1;
defparam ram_block3a61.port_a_first_address = 0;
defparam ram_block3a61.port_a_first_bit_number = 29;
defparam ram_block3a61.port_a_last_address = 8191;
defparam ram_block3a61.port_a_logical_ram_depth = 16384;
defparam ram_block3a61.port_a_logical_ram_width = 32;
defparam ram_block3a61.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_address_clear = "none";
defparam ram_block3a61.port_b_address_clock = "clock1";
defparam ram_block3a61.port_b_address_width = 13;
defparam ram_block3a61.port_b_data_in_clock = "clock1";
defparam ram_block3a61.port_b_data_out_clear = "none";
defparam ram_block3a61.port_b_data_out_clock = "none";
defparam ram_block3a61.port_b_data_width = 1;
defparam ram_block3a61.port_b_first_address = 0;
defparam ram_block3a61.port_b_first_bit_number = 29;
defparam ram_block3a61.port_b_last_address = 8191;
defparam ram_block3a61.port_b_logical_ram_depth = 16384;
defparam ram_block3a61.port_b_logical_ram_width = 32;
defparam ram_block3a61.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a61.port_b_read_enable_clock = "clock1";
defparam ram_block3a61.port_b_write_enable_clock = "clock1";
defparam ram_block3a61.ram_block_type = "M9K";
defparam ram_block3a61.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a61.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X37_Y31_N0
cycloneive_ram_block ram_block3a29(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[29]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[29]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a29_PORTADATAOUT_bus),
	.portbdataout(ram_block3a29_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a29.clk0_core_clock_enable = "ena0";
defparam ram_block3a29.clk1_core_clock_enable = "ena1";
defparam ram_block3a29.data_interleave_offset_in_bits = 1;
defparam ram_block3a29.data_interleave_width_in_bits = 1;
defparam ram_block3a29.init_file = "meminit.hex";
defparam ram_block3a29.init_file_layout = "port_a";
defparam ram_block3a29.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a29.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a29.operation_mode = "bidir_dual_port";
defparam ram_block3a29.port_a_address_clear = "none";
defparam ram_block3a29.port_a_address_width = 13;
defparam ram_block3a29.port_a_byte_enable_clock = "none";
defparam ram_block3a29.port_a_data_out_clear = "none";
defparam ram_block3a29.port_a_data_out_clock = "none";
defparam ram_block3a29.port_a_data_width = 1;
defparam ram_block3a29.port_a_first_address = 0;
defparam ram_block3a29.port_a_first_bit_number = 29;
defparam ram_block3a29.port_a_last_address = 8191;
defparam ram_block3a29.port_a_logical_ram_depth = 16384;
defparam ram_block3a29.port_a_logical_ram_width = 32;
defparam ram_block3a29.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_address_clear = "none";
defparam ram_block3a29.port_b_address_clock = "clock1";
defparam ram_block3a29.port_b_address_width = 13;
defparam ram_block3a29.port_b_data_in_clock = "clock1";
defparam ram_block3a29.port_b_data_out_clear = "none";
defparam ram_block3a29.port_b_data_out_clock = "none";
defparam ram_block3a29.port_b_data_width = 1;
defparam ram_block3a29.port_b_first_address = 0;
defparam ram_block3a29.port_b_first_bit_number = 29;
defparam ram_block3a29.port_b_last_address = 8191;
defparam ram_block3a29.port_b_logical_ram_depth = 16384;
defparam ram_block3a29.port_b_logical_ram_width = 32;
defparam ram_block3a29.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a29.port_b_read_enable_clock = "clock1";
defparam ram_block3a29.port_b_write_enable_clock = "clock1";
defparam ram_block3a29.ram_block_type = "M9K";
defparam ram_block3a29.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a29.mem_init0 = 2048'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000078F3DE001B007700807;
// synopsys translate_on

// Location: M9K_X64_Y28_N0
cycloneive_ram_block ram_block3a62(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a62_PORTADATAOUT_bus),
	.portbdataout(ram_block3a62_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a62.clk0_core_clock_enable = "ena0";
defparam ram_block3a62.clk1_core_clock_enable = "ena1";
defparam ram_block3a62.data_interleave_offset_in_bits = 1;
defparam ram_block3a62.data_interleave_width_in_bits = 1;
defparam ram_block3a62.init_file = "meminit.hex";
defparam ram_block3a62.init_file_layout = "port_a";
defparam ram_block3a62.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a62.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a62.operation_mode = "bidir_dual_port";
defparam ram_block3a62.port_a_address_clear = "none";
defparam ram_block3a62.port_a_address_width = 13;
defparam ram_block3a62.port_a_byte_enable_clock = "none";
defparam ram_block3a62.port_a_data_out_clear = "none";
defparam ram_block3a62.port_a_data_out_clock = "none";
defparam ram_block3a62.port_a_data_width = 1;
defparam ram_block3a62.port_a_first_address = 0;
defparam ram_block3a62.port_a_first_bit_number = 30;
defparam ram_block3a62.port_a_last_address = 8191;
defparam ram_block3a62.port_a_logical_ram_depth = 16384;
defparam ram_block3a62.port_a_logical_ram_width = 32;
defparam ram_block3a62.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_address_clear = "none";
defparam ram_block3a62.port_b_address_clock = "clock1";
defparam ram_block3a62.port_b_address_width = 13;
defparam ram_block3a62.port_b_data_in_clock = "clock1";
defparam ram_block3a62.port_b_data_out_clear = "none";
defparam ram_block3a62.port_b_data_out_clock = "none";
defparam ram_block3a62.port_b_data_width = 1;
defparam ram_block3a62.port_b_first_address = 0;
defparam ram_block3a62.port_b_first_bit_number = 30;
defparam ram_block3a62.port_b_last_address = 8191;
defparam ram_block3a62.port_b_logical_ram_depth = 16384;
defparam ram_block3a62.port_b_logical_ram_width = 32;
defparam ram_block3a62.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a62.port_b_read_enable_clock = "clock1";
defparam ram_block3a62.port_b_write_enable_clock = "clock1";
defparam ram_block3a62.ram_block_type = "M9K";
defparam ram_block3a62.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a62.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X51_Y28_N0
cycloneive_ram_block ram_block3a30(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[30]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[30]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a30_PORTADATAOUT_bus),
	.portbdataout(ram_block3a30_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a30.clk0_core_clock_enable = "ena0";
defparam ram_block3a30.clk1_core_clock_enable = "ena1";
defparam ram_block3a30.data_interleave_offset_in_bits = 1;
defparam ram_block3a30.data_interleave_width_in_bits = 1;
defparam ram_block3a30.init_file = "meminit.hex";
defparam ram_block3a30.init_file_layout = "port_a";
defparam ram_block3a30.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a30.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a30.operation_mode = "bidir_dual_port";
defparam ram_block3a30.port_a_address_clear = "none";
defparam ram_block3a30.port_a_address_width = 13;
defparam ram_block3a30.port_a_byte_enable_clock = "none";
defparam ram_block3a30.port_a_data_out_clear = "none";
defparam ram_block3a30.port_a_data_out_clock = "none";
defparam ram_block3a30.port_a_data_width = 1;
defparam ram_block3a30.port_a_first_address = 0;
defparam ram_block3a30.port_a_first_bit_number = 30;
defparam ram_block3a30.port_a_last_address = 8191;
defparam ram_block3a30.port_a_logical_ram_depth = 16384;
defparam ram_block3a30.port_a_logical_ram_width = 32;
defparam ram_block3a30.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_address_clear = "none";
defparam ram_block3a30.port_b_address_clock = "clock1";
defparam ram_block3a30.port_b_address_width = 13;
defparam ram_block3a30.port_b_data_in_clock = "clock1";
defparam ram_block3a30.port_b_data_out_clear = "none";
defparam ram_block3a30.port_b_data_out_clock = "none";
defparam ram_block3a30.port_b_data_width = 1;
defparam ram_block3a30.port_b_first_address = 0;
defparam ram_block3a30.port_b_first_bit_number = 30;
defparam ram_block3a30.port_b_last_address = 8191;
defparam ram_block3a30.port_b_logical_ram_depth = 16384;
defparam ram_block3a30.port_b_logical_ram_width = 32;
defparam ram_block3a30.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a30.port_b_read_enable_clock = "clock1";
defparam ram_block3a30.port_b_write_enable_clock = "clock1";
defparam ram_block3a30.ram_block_type = "M9K";
defparam ram_block3a30.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a30.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000002000000;
// synopsys translate_on

// Location: M9K_X64_Y22_N0
cycloneive_ram_block ram_block3a63(
	.portawe(\decode4|eq_node[1]~0_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[1]~0_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(!ramaddr),
	.ena1(ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a63_PORTADATAOUT_bus),
	.portbdataout(ram_block3a63_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a63.clk0_core_clock_enable = "ena0";
defparam ram_block3a63.clk1_core_clock_enable = "ena1";
defparam ram_block3a63.data_interleave_offset_in_bits = 1;
defparam ram_block3a63.data_interleave_width_in_bits = 1;
defparam ram_block3a63.init_file = "meminit.hex";
defparam ram_block3a63.init_file_layout = "port_a";
defparam ram_block3a63.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a63.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a63.operation_mode = "bidir_dual_port";
defparam ram_block3a63.port_a_address_clear = "none";
defparam ram_block3a63.port_a_address_width = 13;
defparam ram_block3a63.port_a_byte_enable_clock = "none";
defparam ram_block3a63.port_a_data_out_clear = "none";
defparam ram_block3a63.port_a_data_out_clock = "none";
defparam ram_block3a63.port_a_data_width = 1;
defparam ram_block3a63.port_a_first_address = 0;
defparam ram_block3a63.port_a_first_bit_number = 31;
defparam ram_block3a63.port_a_last_address = 8191;
defparam ram_block3a63.port_a_logical_ram_depth = 16384;
defparam ram_block3a63.port_a_logical_ram_width = 32;
defparam ram_block3a63.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_address_clear = "none";
defparam ram_block3a63.port_b_address_clock = "clock1";
defparam ram_block3a63.port_b_address_width = 13;
defparam ram_block3a63.port_b_data_in_clock = "clock1";
defparam ram_block3a63.port_b_data_out_clear = "none";
defparam ram_block3a63.port_b_data_out_clock = "none";
defparam ram_block3a63.port_b_data_width = 1;
defparam ram_block3a63.port_b_first_address = 0;
defparam ram_block3a63.port_b_first_bit_number = 31;
defparam ram_block3a63.port_b_last_address = 8191;
defparam ram_block3a63.port_b_logical_ram_depth = 16384;
defparam ram_block3a63.port_b_logical_ram_width = 32;
defparam ram_block3a63.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a63.port_b_read_enable_clock = "clock1";
defparam ram_block3a63.port_b_write_enable_clock = "clock1";
defparam ram_block3a63.ram_block_type = "M9K";
defparam ram_block3a63.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a63.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
// synopsys translate_on

// Location: M9K_X64_Y21_N0
cycloneive_ram_block ram_block3a31(
	.portawe(\decode4|eq_node[0]~1_combout ),
	.portare(vcc),
	.portaaddrstall(gnd),
	.portbwe(\decode5|eq_node[0]~1_combout ),
	.portbre(vcc),
	.portbaddrstall(gnd),
	.clk0(clock0),
	.clk1(clock1),
	.ena0(ramaddr),
	.ena1(!ram_rom_addr_reg_13),
	.ena2(vcc),
	.ena3(vcc),
	.clr0(gnd),
	.clr1(gnd),
	.portadatain({data_a[31]}),
	.portaaddr({address_a[12],address_a[11],address_a[10],address_a[9],address_a[8],address_a[7],address_a[6],address_a[5],address_a[4],address_a[3],address_a[2],address_a[1],address_a[0]}),
	.portabyteenamasks(1'b1),
	.portbdatain({data_b[31]}),
	.portbaddr({address_b[12],address_b[11],address_b[10],address_b[9],address_b[8],address_b[7],address_b[6],address_b[5],address_b[4],address_b[3],address_b[2],address_b[1],address_b[0]}),
	.portbbyteenamasks(1'b1),
	.devclrn(devclrn),
	.devpor(devpor),
	.portadataout(ram_block3a31_PORTADATAOUT_bus),
	.portbdataout(ram_block3a31_PORTBDATAOUT_bus));
// synopsys translate_off
defparam ram_block3a31.clk0_core_clock_enable = "ena0";
defparam ram_block3a31.clk1_core_clock_enable = "ena1";
defparam ram_block3a31.data_interleave_offset_in_bits = 1;
defparam ram_block3a31.data_interleave_width_in_bits = 1;
defparam ram_block3a31.init_file = "meminit.hex";
defparam ram_block3a31.init_file_layout = "port_a";
defparam ram_block3a31.logical_ram_name = "ram:RAM|altsyncram:altsyncram_component|altsyncram_99f1:auto_generated|altsyncram_fta2:altsyncram1|ALTSYNCRAM";
defparam ram_block3a31.mixed_port_feed_through_mode = "dont_care";
defparam ram_block3a31.operation_mode = "bidir_dual_port";
defparam ram_block3a31.port_a_address_clear = "none";
defparam ram_block3a31.port_a_address_width = 13;
defparam ram_block3a31.port_a_byte_enable_clock = "none";
defparam ram_block3a31.port_a_data_out_clear = "none";
defparam ram_block3a31.port_a_data_out_clock = "none";
defparam ram_block3a31.port_a_data_width = 1;
defparam ram_block3a31.port_a_first_address = 0;
defparam ram_block3a31.port_a_first_bit_number = 31;
defparam ram_block3a31.port_a_last_address = 8191;
defparam ram_block3a31.port_a_logical_ram_depth = 16384;
defparam ram_block3a31.port_a_logical_ram_width = 32;
defparam ram_block3a31.port_a_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_address_clear = "none";
defparam ram_block3a31.port_b_address_clock = "clock1";
defparam ram_block3a31.port_b_address_width = 13;
defparam ram_block3a31.port_b_data_in_clock = "clock1";
defparam ram_block3a31.port_b_data_out_clear = "none";
defparam ram_block3a31.port_b_data_out_clock = "none";
defparam ram_block3a31.port_b_data_width = 1;
defparam ram_block3a31.port_b_first_address = 0;
defparam ram_block3a31.port_b_first_bit_number = 31;
defparam ram_block3a31.port_b_last_address = 8191;
defparam ram_block3a31.port_b_logical_ram_depth = 16384;
defparam ram_block3a31.port_b_logical_ram_width = 32;
defparam ram_block3a31.port_b_read_during_write_mode = "new_data_with_nbe_read";
defparam ram_block3a31.port_b_read_enable_clock = "clock1";
defparam ram_block3a31.port_b_write_enable_clock = "clock1";
defparam ram_block3a31.ram_block_type = "M9K";
defparam ram_block3a31.mem_init3 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init2 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init1 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
defparam ram_block3a31.mem_init0 = 2048'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000C18426089282400008;
// synopsys translate_on

// Location: FF_X59_Y29_N17
dffeas \address_reg_a[0] (
	.clk(clock0),
	.d(gnd),
	.asdata(ramaddr1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_a_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_a[0] .is_wysiwyg = "true";
defparam \address_reg_a[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N13
dffeas \address_reg_b[0] (
	.clk(clock1),
	.d(\address_reg_b[0]~feeder_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(address_reg_b_0),
	.prn(vcc));
// synopsys translate_off
defparam \address_reg_b[0] .is_wysiwyg = "true";
defparam \address_reg_b[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N12
cycloneive_lcell_comb \address_reg_b[0]~feeder (
// Equation(s):
// \address_reg_b[0]~feeder_combout  = ram_rom_addr_reg_13

	.dataa(gnd),
	.datab(gnd),
	.datac(ram_rom_addr_reg_13),
	.datad(gnd),
	.cin(gnd),
	.combout(\address_reg_b[0]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \address_reg_b[0]~feeder .lut_mask = 16'hF0F0;
defparam \address_reg_b[0]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa (
	ramaddr,
	ramWEN,
	always1,
	eq_node_1,
	eq_node_0,
	devpor,
	devclrn,
	devoe);
input 	ramaddr;
input 	ramWEN;
input 	always1;
output 	eq_node_1;
output 	eq_node_0;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X59_Y29_N24
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (!\ramWEN~0_combout  & (!\ramaddr~29_combout  & always1))

	.dataa(ramWEN),
	.datab(gnd),
	.datac(ramaddr),
	.datad(always1),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h0500;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X59_Y29_N22
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (!\ramWEN~0_combout  & (\ramaddr~29_combout  & always1))

	.dataa(ramWEN),
	.datab(gnd),
	.datac(ramaddr),
	.datad(always1),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h5000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module decode_jsa_1 (
	ram_rom_addr_reg_13,
	sdr,
	eq_node_1,
	eq_node_0,
	irf_reg_2_1,
	state_5,
	devpor,
	devclrn,
	devoe);
input 	ram_rom_addr_reg_13;
input 	sdr;
output 	eq_node_1;
output 	eq_node_0;
input 	irf_reg_2_1;
input 	state_5;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;



// Location: LCCOMB_X46_Y32_N18
cycloneive_lcell_comb \eq_node[1]~0 (
// Equation(s):
// eq_node_1 = (ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & sdr)))

	.dataa(ram_rom_addr_reg_13),
	.datab(irf_reg_2_1),
	.datac(state_5),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_1),
	.cout());
// synopsys translate_off
defparam \eq_node[1]~0 .lut_mask = 16'h8000;
defparam \eq_node[1]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N4
cycloneive_lcell_comb \eq_node[0]~1 (
// Equation(s):
// eq_node_0 = (!ram_rom_addr_reg_13 & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|irf_reg[1][2]~q  & (\auto_hub|jtag_hub_gen:sld_jtag_hub_inst|shadow_jsm|state [5] & sdr)))

	.dataa(ram_rom_addr_reg_13),
	.datab(irf_reg_2_1),
	.datac(state_5),
	.datad(sdr),
	.cin(gnd),
	.combout(eq_node_0),
	.cout());
// synopsys translate_off
defparam \eq_node[0]~1 .lut_mask = 16'h4000;
defparam \eq_node[0]~1 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_mod_ram_rom (
	ram_block3a32,
	ram_block3a0,
	ram_block3a33,
	ram_block3a1,
	ram_block3a34,
	ram_block3a2,
	ram_block3a35,
	ram_block3a3,
	ram_block3a36,
	ram_block3a4,
	ram_block3a37,
	ram_block3a5,
	ram_block3a38,
	ram_block3a6,
	ram_block3a39,
	ram_block3a7,
	ram_block3a40,
	ram_block3a8,
	ram_block3a41,
	ram_block3a9,
	ram_block3a42,
	ram_block3a10,
	ram_block3a43,
	ram_block3a11,
	ram_block3a44,
	ram_block3a12,
	ram_block3a45,
	ram_block3a13,
	ram_block3a46,
	ram_block3a14,
	ram_block3a47,
	ram_block3a15,
	ram_block3a48,
	ram_block3a16,
	ram_block3a49,
	ram_block3a17,
	ram_block3a50,
	ram_block3a18,
	ram_block3a51,
	ram_block3a19,
	ram_block3a52,
	ram_block3a20,
	ram_block3a53,
	ram_block3a21,
	ram_block3a54,
	ram_block3a22,
	ram_block3a55,
	ram_block3a23,
	ram_block3a56,
	ram_block3a24,
	ram_block3a57,
	ram_block3a25,
	ram_block3a58,
	ram_block3a26,
	ram_block3a59,
	ram_block3a27,
	ram_block3a60,
	ram_block3a28,
	ram_block3a61,
	ram_block3a29,
	ram_block3a62,
	ram_block3a30,
	ram_block3a63,
	ram_block3a31,
	is_in_use_reg1,
	ram_rom_data_reg_0,
	ram_rom_addr_reg_13,
	ram_rom_addr_reg_0,
	ram_rom_addr_reg_1,
	ram_rom_addr_reg_2,
	ram_rom_addr_reg_3,
	ram_rom_addr_reg_4,
	ram_rom_addr_reg_5,
	ram_rom_addr_reg_6,
	ram_rom_addr_reg_7,
	ram_rom_addr_reg_8,
	ram_rom_addr_reg_9,
	ram_rom_addr_reg_10,
	ram_rom_addr_reg_11,
	ram_rom_addr_reg_12,
	ram_rom_data_reg_1,
	ram_rom_data_reg_2,
	ram_rom_data_reg_3,
	ram_rom_data_reg_4,
	ram_rom_data_reg_5,
	ram_rom_data_reg_6,
	ram_rom_data_reg_7,
	ram_rom_data_reg_8,
	ram_rom_data_reg_9,
	ram_rom_data_reg_10,
	ram_rom_data_reg_11,
	ram_rom_data_reg_12,
	ram_rom_data_reg_13,
	ram_rom_data_reg_14,
	ram_rom_data_reg_15,
	ram_rom_data_reg_16,
	ram_rom_data_reg_17,
	ram_rom_data_reg_18,
	ram_rom_data_reg_19,
	ram_rom_data_reg_20,
	ram_rom_data_reg_21,
	ram_rom_data_reg_22,
	ram_rom_data_reg_23,
	ram_rom_data_reg_24,
	ram_rom_data_reg_25,
	ram_rom_data_reg_26,
	ram_rom_data_reg_27,
	ram_rom_data_reg_28,
	ram_rom_data_reg_29,
	ram_rom_data_reg_30,
	ram_rom_data_reg_31,
	ir_loaded_address_reg_0,
	ir_loaded_address_reg_1,
	ir_loaded_address_reg_2,
	ir_loaded_address_reg_3,
	tdo,
	sdr,
	address_reg_b_0,
	altera_internal_jtag,
	state_4,
	ir_in,
	irf_reg_1_1,
	irf_reg_2_1,
	irf_reg_4_1,
	node_ena_1,
	clr,
	virtual_ir_scan_reg,
	state_3,
	state_5,
	state_8,
	raw_tck,
	devpor,
	devclrn,
	devoe);
input 	ram_block3a32;
input 	ram_block3a0;
input 	ram_block3a33;
input 	ram_block3a1;
input 	ram_block3a34;
input 	ram_block3a2;
input 	ram_block3a35;
input 	ram_block3a3;
input 	ram_block3a36;
input 	ram_block3a4;
input 	ram_block3a37;
input 	ram_block3a5;
input 	ram_block3a38;
input 	ram_block3a6;
input 	ram_block3a39;
input 	ram_block3a7;
input 	ram_block3a40;
input 	ram_block3a8;
input 	ram_block3a41;
input 	ram_block3a9;
input 	ram_block3a42;
input 	ram_block3a10;
input 	ram_block3a43;
input 	ram_block3a11;
input 	ram_block3a44;
input 	ram_block3a12;
input 	ram_block3a45;
input 	ram_block3a13;
input 	ram_block3a46;
input 	ram_block3a14;
input 	ram_block3a47;
input 	ram_block3a15;
input 	ram_block3a48;
input 	ram_block3a16;
input 	ram_block3a49;
input 	ram_block3a17;
input 	ram_block3a50;
input 	ram_block3a18;
input 	ram_block3a51;
input 	ram_block3a19;
input 	ram_block3a52;
input 	ram_block3a20;
input 	ram_block3a53;
input 	ram_block3a21;
input 	ram_block3a54;
input 	ram_block3a22;
input 	ram_block3a55;
input 	ram_block3a23;
input 	ram_block3a56;
input 	ram_block3a24;
input 	ram_block3a57;
input 	ram_block3a25;
input 	ram_block3a58;
input 	ram_block3a26;
input 	ram_block3a59;
input 	ram_block3a27;
input 	ram_block3a60;
input 	ram_block3a28;
input 	ram_block3a61;
input 	ram_block3a29;
input 	ram_block3a62;
input 	ram_block3a30;
input 	ram_block3a63;
input 	ram_block3a31;
output 	is_in_use_reg1;
output 	ram_rom_data_reg_0;
output 	ram_rom_addr_reg_13;
output 	ram_rom_addr_reg_0;
output 	ram_rom_addr_reg_1;
output 	ram_rom_addr_reg_2;
output 	ram_rom_addr_reg_3;
output 	ram_rom_addr_reg_4;
output 	ram_rom_addr_reg_5;
output 	ram_rom_addr_reg_6;
output 	ram_rom_addr_reg_7;
output 	ram_rom_addr_reg_8;
output 	ram_rom_addr_reg_9;
output 	ram_rom_addr_reg_10;
output 	ram_rom_addr_reg_11;
output 	ram_rom_addr_reg_12;
output 	ram_rom_data_reg_1;
output 	ram_rom_data_reg_2;
output 	ram_rom_data_reg_3;
output 	ram_rom_data_reg_4;
output 	ram_rom_data_reg_5;
output 	ram_rom_data_reg_6;
output 	ram_rom_data_reg_7;
output 	ram_rom_data_reg_8;
output 	ram_rom_data_reg_9;
output 	ram_rom_data_reg_10;
output 	ram_rom_data_reg_11;
output 	ram_rom_data_reg_12;
output 	ram_rom_data_reg_13;
output 	ram_rom_data_reg_14;
output 	ram_rom_data_reg_15;
output 	ram_rom_data_reg_16;
output 	ram_rom_data_reg_17;
output 	ram_rom_data_reg_18;
output 	ram_rom_data_reg_19;
output 	ram_rom_data_reg_20;
output 	ram_rom_data_reg_21;
output 	ram_rom_data_reg_22;
output 	ram_rom_data_reg_23;
output 	ram_rom_data_reg_24;
output 	ram_rom_data_reg_25;
output 	ram_rom_data_reg_26;
output 	ram_rom_data_reg_27;
output 	ram_rom_data_reg_28;
output 	ram_rom_data_reg_29;
output 	ram_rom_data_reg_30;
output 	ram_rom_data_reg_31;
output 	ir_loaded_address_reg_0;
output 	ir_loaded_address_reg_1;
output 	ir_loaded_address_reg_2;
output 	ir_loaded_address_reg_3;
output 	tdo;
output 	sdr;
input 	address_reg_b_0;
input 	altera_internal_jtag;
input 	state_4;
input 	[4:0] ir_in;
input 	irf_reg_1_1;
input 	irf_reg_2_1;
input 	irf_reg_4_1;
input 	node_ena_1;
input 	clr;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_5;
input 	state_8;
input 	raw_tck;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \Add1~1 ;
wire \Add1~0_combout ;
wire \Add1~3 ;
wire \Add1~2_combout ;
wire \Add1~5 ;
wire \Add1~4_combout ;
wire \Add1~7 ;
wire \Add1~6_combout ;
wire \Add1~9 ;
wire \Add1~8_combout ;
wire \Add1~10_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~8_combout ;
wire \is_in_use_reg~0_combout ;
wire \ram_rom_data_reg[0]~0_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~4_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~12_combout ;
wire \ram_rom_data_shift_cntr_reg[3]~11_combout ;
wire \ram_rom_data_shift_cntr_reg[2]~9_combout ;
wire \ram_rom_data_shift_cntr_reg[5]~10_combout ;
wire \ram_rom_data_shift_cntr_reg[4]~7_combout ;
wire \Equal1~0_combout ;
wire \ram_rom_data_shift_cntr_reg[0]~6_combout ;
wire \Equal1~1_combout ;
wire \ram_rom_data_shift_cntr_reg[1]~5_combout ;
wire \process_0~2_combout ;
wire \ram_rom_data_reg[9]~32_combout ;
wire \ram_rom_addr_reg[0]~15 ;
wire \ram_rom_addr_reg[1]~17 ;
wire \ram_rom_addr_reg[2]~19 ;
wire \ram_rom_addr_reg[3]~21 ;
wire \ram_rom_addr_reg[4]~23 ;
wire \ram_rom_addr_reg[5]~25 ;
wire \ram_rom_addr_reg[6]~27 ;
wire \ram_rom_addr_reg[7]~29 ;
wire \ram_rom_addr_reg[8]~31 ;
wire \ram_rom_addr_reg[9]~33 ;
wire \ram_rom_addr_reg[10]~35 ;
wire \ram_rom_addr_reg[11]~37 ;
wire \ram_rom_addr_reg[12]~39 ;
wire \ram_rom_addr_reg[13]~40_combout ;
wire \process_0~3_combout ;
wire \ram_rom_addr_reg[7]~42_combout ;
wire \ram_rom_addr_reg[7]~43_combout ;
wire \ram_rom_addr_reg[0]~14_combout ;
wire \ram_rom_addr_reg[1]~16_combout ;
wire \ram_rom_addr_reg[2]~18_combout ;
wire \ram_rom_addr_reg[3]~20_combout ;
wire \ram_rom_addr_reg[4]~22_combout ;
wire \ram_rom_addr_reg[5]~24_combout ;
wire \ram_rom_addr_reg[6]~26_combout ;
wire \ram_rom_addr_reg[7]~28_combout ;
wire \ram_rom_addr_reg[8]~30_combout ;
wire \ram_rom_addr_reg[9]~32_combout ;
wire \ram_rom_addr_reg[10]~34_combout ;
wire \ram_rom_addr_reg[11]~36_combout ;
wire \ram_rom_addr_reg[12]~38_combout ;
wire \ram_rom_data_reg[1]~1_combout ;
wire \ram_rom_data_reg[2]~2_combout ;
wire \ram_rom_data_reg[3]~3_combout ;
wire \ram_rom_data_reg[4]~4_combout ;
wire \ram_rom_data_reg[5]~5_combout ;
wire \ram_rom_data_reg[6]~6_combout ;
wire \ram_rom_data_reg[7]~7_combout ;
wire \ram_rom_data_reg[8]~8_combout ;
wire \ram_rom_data_reg[9]~9_combout ;
wire \ram_rom_data_reg[10]~10_combout ;
wire \ram_rom_data_reg[11]~11_combout ;
wire \ram_rom_data_reg[12]~12_combout ;
wire \ram_rom_data_reg[13]~13_combout ;
wire \ram_rom_data_reg[14]~14_combout ;
wire \ram_rom_data_reg[15]~15_combout ;
wire \ram_rom_data_reg[16]~16_combout ;
wire \ram_rom_data_reg[17]~17_combout ;
wire \ram_rom_data_reg[18]~18_combout ;
wire \ram_rom_data_reg[19]~19_combout ;
wire \ram_rom_data_reg[20]~20_combout ;
wire \ram_rom_data_reg[21]~21_combout ;
wire \ram_rom_data_reg[22]~22_combout ;
wire \ram_rom_data_reg[23]~23_combout ;
wire \ram_rom_data_reg[24]~24_combout ;
wire \ram_rom_data_reg[25]~25_combout ;
wire \ram_rom_data_reg[26]~26_combout ;
wire \ram_rom_data_reg[27]~27_combout ;
wire \ram_rom_data_reg[28]~28_combout ;
wire \ram_rom_data_reg[29]~29_combout ;
wire \ram_rom_data_reg[30]~30_combout ;
wire \ram_rom_data_reg[31]~31_combout ;
wire \process_0~0_combout ;
wire \process_0~1_combout ;
wire \ir_loaded_address_reg[1]~feeder_combout ;
wire \ir_loaded_address_reg[2]~feeder_combout ;
wire \bypass_reg_out~0_combout ;
wire \bypass_reg_out~q ;
wire \tdo~0_combout ;
wire [5:0] ram_rom_data_shift_cntr_reg;
wire [3:0] \ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR ;


sld_rom_sr \ram_rom_logic_gen:name_gen:info_rom_sr (
	.WORD_SR_0(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.sdr(sdr),
	.altera_internal_jtag(altera_internal_jtag),
	.state_4(state_4),
	.virtual_ir_scan_reg(virtual_ir_scan_reg),
	.state_3(state_3),
	.state_8(state_8),
	.TCK(raw_tck),
	.devpor(devpor),
	.devclrn(devclrn),
	.devoe(devoe));

// Location: LCCOMB_X45_Y32_N4
cycloneive_lcell_comb \Add1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\Add1~0_combout ),
	.cout(\Add1~1 ));
// synopsys translate_off
defparam \Add1~0 .lut_mask = 16'h55AA;
defparam \Add1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N6
cycloneive_lcell_comb \Add1~2 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~1 ),
	.combout(\Add1~2_combout ),
	.cout(\Add1~3 ));
// synopsys translate_off
defparam \Add1~2 .lut_mask = 16'h3C3F;
defparam \Add1~2 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N8
cycloneive_lcell_comb \Add1~4 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~3 ),
	.combout(\Add1~4_combout ),
	.cout(\Add1~5 ));
// synopsys translate_off
defparam \Add1~4 .lut_mask = 16'hC30C;
defparam \Add1~4 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N10
cycloneive_lcell_comb \Add1~6 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~5 ),
	.combout(\Add1~6_combout ),
	.cout(\Add1~7 ));
// synopsys translate_off
defparam \Add1~6 .lut_mask = 16'h5A5F;
defparam \Add1~6 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N12
cycloneive_lcell_comb \Add1~8 (
	.dataa(gnd),
	.datab(ram_rom_data_shift_cntr_reg[4]),
	.datac(gnd),
	.datad(vcc),
	.cin(\Add1~7 ),
	.combout(\Add1~8_combout ),
	.cout(\Add1~9 ));
// synopsys translate_off
defparam \Add1~8 .lut_mask = 16'hC30C;
defparam \Add1~8 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N14
cycloneive_lcell_comb \Add1~10 (
	.dataa(ram_rom_data_shift_cntr_reg[5]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.cin(\Add1~9 ),
	.combout(\Add1~10_combout ),
	.cout());
// synopsys translate_off
defparam \Add1~10 .lut_mask = 16'h5A5A;
defparam \Add1~10 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X45_Y32_N31
dffeas \ram_rom_data_shift_cntr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[3]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N30
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~8 (
	.dataa(\Add1~6_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datac(ram_rom_data_shift_cntr_reg[3]),
	.datad(\ram_rom_data_shift_cntr_reg[3]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~8 .lut_mask = 16'hF222;
defparam \ram_rom_data_shift_cntr_reg[3]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X48_Y32_N5
dffeas is_in_use_reg(
	.clk(raw_tck),
	.d(\is_in_use_reg~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(ir_in[0]),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(is_in_use_reg1),
	.prn(vcc));
// synopsys translate_off
defparam is_in_use_reg.is_wysiwyg = "true";
defparam is_in_use_reg.power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N21
dffeas \ram_rom_data_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[0]~0_combout ),
	.asdata(ram_rom_data_reg_1),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N29
dffeas \ram_rom_addr_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[13]~40_combout ),
	.asdata(altera_internal_jtag),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N3
dffeas \ram_rom_addr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[0]~14_combout ),
	.asdata(ram_rom_addr_reg_1),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N5
dffeas \ram_rom_addr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[1]~16_combout ),
	.asdata(ram_rom_addr_reg_2),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N7
dffeas \ram_rom_addr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[2]~18_combout ),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N9
dffeas \ram_rom_addr_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[3]~20_combout ),
	.asdata(ram_rom_addr_reg_4),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N11
dffeas \ram_rom_addr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[4]~22_combout ),
	.asdata(ram_rom_addr_reg_5),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N13
dffeas \ram_rom_addr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[5]~24_combout ),
	.asdata(ram_rom_addr_reg_6),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N15
dffeas \ram_rom_addr_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[6]~26_combout ),
	.asdata(ram_rom_addr_reg_7),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N17
dffeas \ram_rom_addr_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[7]~28_combout ),
	.asdata(ram_rom_addr_reg_8),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N19
dffeas \ram_rom_addr_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[8]~30_combout ),
	.asdata(ram_rom_addr_reg_9),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N21
dffeas \ram_rom_addr_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[9]~32_combout ),
	.asdata(ram_rom_addr_reg_10),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N23
dffeas \ram_rom_addr_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[10]~34_combout ),
	.asdata(ram_rom_addr_reg_11),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N25
dffeas \ram_rom_addr_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[11]~36_combout ),
	.asdata(ram_rom_addr_reg_12),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X49_Y32_N27
dffeas \ram_rom_addr_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_addr_reg[12]~38_combout ),
	.asdata(ram_rom_addr_reg_13),
	.clrn(!ir_in[0]),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~3_combout ),
	.ena(\ram_rom_addr_reg[7]~43_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_addr_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_addr_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_addr_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N15
dffeas \ram_rom_data_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[1]~1_combout ),
	.asdata(ram_rom_data_reg_2),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N9
dffeas \ram_rom_data_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[2]~2_combout ),
	.asdata(ram_rom_data_reg_3),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N23
dffeas \ram_rom_data_reg[3] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[3]~3_combout ),
	.asdata(ram_rom_data_reg_4),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[3] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[3] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N25
dffeas \ram_rom_data_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[4]~4_combout ),
	.asdata(ram_rom_data_reg_5),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_4),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[4] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N25
dffeas \ram_rom_data_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[5]~5_combout ),
	.asdata(ram_rom_data_reg_6),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_5),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[5] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N19
dffeas \ram_rom_data_reg[6] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[6]~6_combout ),
	.asdata(ram_rom_data_reg_7),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_6),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[6] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[6] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N21
dffeas \ram_rom_data_reg[7] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[7]~7_combout ),
	.asdata(ram_rom_data_reg_8),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_7),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[7] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[7] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N31
dffeas \ram_rom_data_reg[8] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[8]~8_combout ),
	.asdata(ram_rom_data_reg_9),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_8),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[8] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[8] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N17
dffeas \ram_rom_data_reg[9] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[9]~9_combout ),
	.asdata(ram_rom_data_reg_10),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_9),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[9] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[9] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N11
dffeas \ram_rom_data_reg[10] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[10]~10_combout ),
	.asdata(ram_rom_data_reg_11),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_10),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[10] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[10] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N29
dffeas \ram_rom_data_reg[11] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[11]~11_combout ),
	.asdata(ram_rom_data_reg_12),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_11),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[11] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[11] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N27
dffeas \ram_rom_data_reg[12] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[12]~12_combout ),
	.asdata(ram_rom_data_reg_13),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_12),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[12] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[12] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N9
dffeas \ram_rom_data_reg[13] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[13]~13_combout ),
	.asdata(ram_rom_data_reg_14),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_13),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[13] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[13] .power_up = "low";
// synopsys translate_on

// Location: FF_X75_Y31_N15
dffeas \ram_rom_data_reg[14] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[14]~14_combout ),
	.asdata(ram_rom_data_reg_15),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_14),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[14] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[14] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N27
dffeas \ram_rom_data_reg[15] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[15]~15_combout ),
	.asdata(ram_rom_data_reg_16),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_15),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[15] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[15] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N29
dffeas \ram_rom_data_reg[16] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[16]~16_combout ),
	.asdata(ram_rom_data_reg_17),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_16),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[16] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[16] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N27
dffeas \ram_rom_data_reg[17] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[17]~17_combout ),
	.asdata(ram_rom_data_reg_18),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_17),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[17] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[17] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N1
dffeas \ram_rom_data_reg[18] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[18]~18_combout ),
	.asdata(ram_rom_data_reg_19),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_18),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[18] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[18] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N23
dffeas \ram_rom_data_reg[19] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[19]~19_combout ),
	.asdata(ram_rom_data_reg_20),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_19),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[19] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[19] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N9
dffeas \ram_rom_data_reg[20] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[20]~20_combout ),
	.asdata(ram_rom_data_reg_21),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_20),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[20] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[20] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N19
dffeas \ram_rom_data_reg[21] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[21]~21_combout ),
	.asdata(ram_rom_data_reg_22),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_21),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[21] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[21] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N5
dffeas \ram_rom_data_reg[22] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[22]~22_combout ),
	.asdata(ram_rom_data_reg_23),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_22),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[22] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[22] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N31
dffeas \ram_rom_data_reg[23] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[23]~23_combout ),
	.asdata(ram_rom_data_reg_24),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_23),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[23] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[23] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N13
dffeas \ram_rom_data_reg[24] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[24]~24_combout ),
	.asdata(ram_rom_data_reg_25),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_24),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[24] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[24] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N15
dffeas \ram_rom_data_reg[25] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[25]~25_combout ),
	.asdata(ram_rom_data_reg_26),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_25),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[25] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[25] .power_up = "low";
// synopsys translate_on

// Location: FF_X52_Y33_N21
dffeas \ram_rom_data_reg[26] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[26]~26_combout ),
	.asdata(ram_rom_data_reg_27),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_26),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[26] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[26] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N13
dffeas \ram_rom_data_reg[27] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[27]~27_combout ),
	.asdata(ram_rom_data_reg_28),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_27),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[27] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[27] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N19
dffeas \ram_rom_data_reg[28] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[28]~28_combout ),
	.asdata(ram_rom_data_reg_29),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_28),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[28] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[28] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N29
dffeas \ram_rom_data_reg[29] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[29]~29_combout ),
	.asdata(ram_rom_data_reg_30),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_29),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[29] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[29] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N31
dffeas \ram_rom_data_reg[30] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[30]~30_combout ),
	.asdata(ram_rom_data_reg_31),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_30),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[30] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[30] .power_up = "low";
// synopsys translate_on

// Location: FF_X50_Y28_N17
dffeas \ram_rom_data_reg[31] (
	.clk(raw_tck),
	.d(\ram_rom_data_reg[31]~31_combout ),
	.asdata(altera_internal_jtag),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(\process_0~2_combout ),
	.ena(\ram_rom_data_reg[9]~32_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_reg_31),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_reg[31] .is_wysiwyg = "true";
defparam \ram_rom_data_reg[31] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N9
dffeas \ir_loaded_address_reg[0] (
	.clk(raw_tck),
	.d(gnd),
	.asdata(ram_rom_addr_reg_0),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_0),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[0] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[0] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N3
dffeas \ir_loaded_address_reg[1] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[1]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_1),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[1] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[1] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N25
dffeas \ir_loaded_address_reg[2] (
	.clk(raw_tck),
	.d(\ir_loaded_address_reg[2]~feeder_combout ),
	.asdata(vcc),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_2),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[2] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[2] .power_up = "low";
// synopsys translate_on

// Location: FF_X46_Y32_N23
dffeas \ir_loaded_address_reg[3] (
	.clk(raw_tck),
	.d(gnd),
	.asdata(ram_rom_addr_reg_3),
	.clrn(!\process_0~0_combout ),
	.aload(gnd),
	.sclr(gnd),
	.sload(vcc),
	.ena(\process_0~1_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ir_loaded_address_reg_3),
	.prn(vcc));
// synopsys translate_off
defparam \ir_loaded_address_reg[3] .is_wysiwyg = "true";
defparam \ir_loaded_address_reg[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N10
cycloneive_lcell_comb \tdo~1 (
	.dataa(\tdo~0_combout ),
	.datab(\ram_rom_logic_gen:name_gen:info_rom_sr|WORD_SR [0]),
	.datac(ir_in[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(tdo),
	.cout());
// synopsys translate_off
defparam \tdo~1 .lut_mask = 16'hCACA;
defparam \tdo~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N16
cycloneive_lcell_comb \sdr~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(virtual_ir_scan_reg),
	.datad(node_ena_1),
	.cin(gnd),
	.combout(sdr),
	.cout());
// synopsys translate_off
defparam \sdr~0 .lut_mask = 16'h0F00;
defparam \sdr~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X48_Y32_N4
cycloneive_lcell_comb \is_in_use_reg~0 (
	.dataa(gnd),
	.datab(gnd),
	.datac(is_in_use_reg1),
	.datad(irf_reg_4_1),
	.cin(gnd),
	.combout(\is_in_use_reg~0_combout ),
	.cout());
// synopsys translate_off
defparam \is_in_use_reg~0 .lut_mask = 16'h00F0;
defparam \is_in_use_reg~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N20
cycloneive_lcell_comb \ram_rom_data_reg[0]~0 (
	.dataa(ram_block3a0),
	.datab(ram_block3a32),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[0]~0_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[0]~0 .lut_mask = 16'hCCAA;
defparam \ram_rom_data_reg[0]~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N6
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~4 (
	.dataa(sdr),
	.datab(irf_reg_2_1),
	.datac(irf_reg_1_1),
	.datad(state_4),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~4 .lut_mask = 16'hA800;
defparam \ram_rom_data_shift_cntr_reg[5]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N18
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~12 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(\Equal1~0_combout ),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~12 .lut_mask = 16'h8F0F;
defparam \ram_rom_data_shift_cntr_reg[5]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N0
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[3]~11 (
	.dataa(ram_rom_data_shift_cntr_reg[0]),
	.datab(\Equal1~0_combout ),
	.datac(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[3]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[3]~11 .lut_mask = 16'h070F;
defparam \ram_rom_data_shift_cntr_reg[3]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N28
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[2]~9 (
	.dataa(\Add1~4_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datac(ram_rom_data_shift_cntr_reg[2]),
	.datad(\ram_rom_data_shift_cntr_reg[3]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2]~9 .lut_mask = 16'hF222;
defparam \ram_rom_data_shift_cntr_reg[2]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N29
dffeas \ram_rom_data_shift_cntr_reg[2] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[2]~9_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[2]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[2] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N26
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[5]~10 (
	.dataa(\Add1~10_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(\ram_rom_data_shift_cntr_reg[3]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5]~10 .lut_mask = 16'hF222;
defparam \ram_rom_data_shift_cntr_reg[5]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N27
dffeas \ram_rom_data_shift_cntr_reg[5] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[5]~10_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[5]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[5] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[5] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N20
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[4]~7 (
	.dataa(\Add1~8_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datac(ram_rom_data_shift_cntr_reg[4]),
	.datad(\ram_rom_data_shift_cntr_reg[3]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4]~7 .lut_mask = 16'hF222;
defparam \ram_rom_data_shift_cntr_reg[4]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N21
dffeas \ram_rom_data_shift_cntr_reg[4] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[4]~7_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[4]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[4] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N16
cycloneive_lcell_comb \Equal1~0 (
	.dataa(ram_rom_data_shift_cntr_reg[3]),
	.datab(ram_rom_data_shift_cntr_reg[2]),
	.datac(ram_rom_data_shift_cntr_reg[5]),
	.datad(ram_rom_data_shift_cntr_reg[4]),
	.cin(gnd),
	.combout(\Equal1~0_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~0 .lut_mask = 16'h0800;
defparam \Equal1~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N22
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[0]~6 (
	.dataa(\Add1~0_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~12_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(\ram_rom_data_shift_cntr_reg[3]~11_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0]~6 .lut_mask = 16'hF222;
defparam \ram_rom_data_shift_cntr_reg[0]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N23
dffeas \ram_rom_data_shift_cntr_reg[0] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[0]~6_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[0]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[0] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N2
cycloneive_lcell_comb \Equal1~1 (
	.dataa(gnd),
	.datab(\Equal1~0_combout ),
	.datac(ram_rom_data_shift_cntr_reg[0]),
	.datad(gnd),
	.cin(gnd),
	.combout(\Equal1~1_combout ),
	.cout());
// synopsys translate_off
defparam \Equal1~1 .lut_mask = 16'hC0C0;
defparam \Equal1~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X45_Y32_N24
cycloneive_lcell_comb \ram_rom_data_shift_cntr_reg[1]~5 (
	.dataa(\Add1~2_combout ),
	.datab(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.datac(ram_rom_data_shift_cntr_reg[1]),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1]~5 .lut_mask = 16'h08B8;
defparam \ram_rom_data_shift_cntr_reg[1]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X45_Y32_N25
dffeas \ram_rom_data_shift_cntr_reg[1] (
	.clk(raw_tck),
	.d(\ram_rom_data_shift_cntr_reg[1]~5_combout ),
	.asdata(vcc),
	.clrn(!ir_in[3]),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(ram_rom_data_shift_cntr_reg[1]),
	.prn(vcc));
// synopsys translate_off
defparam \ram_rom_data_shift_cntr_reg[1] .is_wysiwyg = "true";
defparam \ram_rom_data_shift_cntr_reg[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N12
cycloneive_lcell_comb \process_0~2 (
	.dataa(irf_reg_1_1),
	.datab(ram_rom_data_shift_cntr_reg[1]),
	.datac(ir_in[3]),
	.datad(\Equal1~1_combout ),
	.cin(gnd),
	.combout(\process_0~2_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~2 .lut_mask = 16'h070F;
defparam \process_0~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N10
cycloneive_lcell_comb \ram_rom_data_reg[9]~32 (
	.dataa(gnd),
	.datab(gnd),
	.datac(\process_0~2_combout ),
	.datad(\ram_rom_data_shift_cntr_reg[5]~4_combout ),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~32_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~32 .lut_mask = 16'hFF0F;
defparam \ram_rom_data_reg[9]~32 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N2
cycloneive_lcell_comb \ram_rom_addr_reg[0]~14 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_0),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[0]~14_combout ),
	.cout(\ram_rom_addr_reg[0]~15 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[0]~14 .lut_mask = 16'h33CC;
defparam \ram_rom_addr_reg[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N4
cycloneive_lcell_comb \ram_rom_addr_reg[1]~16 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_1),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[0]~15 ),
	.combout(\ram_rom_addr_reg[1]~16_combout ),
	.cout(\ram_rom_addr_reg[1]~17 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[1]~16 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[1]~16 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N6
cycloneive_lcell_comb \ram_rom_addr_reg[2]~18 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_2),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[1]~17 ),
	.combout(\ram_rom_addr_reg[2]~18_combout ),
	.cout(\ram_rom_addr_reg[2]~19 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[2]~18 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[2]~18 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N8
cycloneive_lcell_comb \ram_rom_addr_reg[3]~20 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_3),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[2]~19 ),
	.combout(\ram_rom_addr_reg[3]~20_combout ),
	.cout(\ram_rom_addr_reg[3]~21 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[3]~20 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[3]~20 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N10
cycloneive_lcell_comb \ram_rom_addr_reg[4]~22 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_4),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[3]~21 ),
	.combout(\ram_rom_addr_reg[4]~22_combout ),
	.cout(\ram_rom_addr_reg[4]~23 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[4]~22 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[4]~22 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N12
cycloneive_lcell_comb \ram_rom_addr_reg[5]~24 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_5),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[4]~23 ),
	.combout(\ram_rom_addr_reg[5]~24_combout ),
	.cout(\ram_rom_addr_reg[5]~25 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[5]~24 .lut_mask = 16'h3C3F;
defparam \ram_rom_addr_reg[5]~24 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N14
cycloneive_lcell_comb \ram_rom_addr_reg[6]~26 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_6),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[5]~25 ),
	.combout(\ram_rom_addr_reg[6]~26_combout ),
	.cout(\ram_rom_addr_reg[6]~27 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[6]~26 .lut_mask = 16'hC30C;
defparam \ram_rom_addr_reg[6]~26 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N16
cycloneive_lcell_comb \ram_rom_addr_reg[7]~28 (
	.dataa(ram_rom_addr_reg_7),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[6]~27 ),
	.combout(\ram_rom_addr_reg[7]~28_combout ),
	.cout(\ram_rom_addr_reg[7]~29 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~28 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[7]~28 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N18
cycloneive_lcell_comb \ram_rom_addr_reg[8]~30 (
	.dataa(ram_rom_addr_reg_8),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[7]~29 ),
	.combout(\ram_rom_addr_reg[8]~30_combout ),
	.cout(\ram_rom_addr_reg[8]~31 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[8]~30 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[8]~30 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N20
cycloneive_lcell_comb \ram_rom_addr_reg[9]~32 (
	.dataa(ram_rom_addr_reg_9),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[8]~31 ),
	.combout(\ram_rom_addr_reg[9]~32_combout ),
	.cout(\ram_rom_addr_reg[9]~33 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[9]~32 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[9]~32 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N22
cycloneive_lcell_comb \ram_rom_addr_reg[10]~34 (
	.dataa(ram_rom_addr_reg_10),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[9]~33 ),
	.combout(\ram_rom_addr_reg[10]~34_combout ),
	.cout(\ram_rom_addr_reg[10]~35 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[10]~34 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[10]~34 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N24
cycloneive_lcell_comb \ram_rom_addr_reg[11]~36 (
	.dataa(ram_rom_addr_reg_11),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[10]~35 ),
	.combout(\ram_rom_addr_reg[11]~36_combout ),
	.cout(\ram_rom_addr_reg[11]~37 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[11]~36 .lut_mask = 16'h5A5F;
defparam \ram_rom_addr_reg[11]~36 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N26
cycloneive_lcell_comb \ram_rom_addr_reg[12]~38 (
	.dataa(ram_rom_addr_reg_12),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\ram_rom_addr_reg[11]~37 ),
	.combout(\ram_rom_addr_reg[12]~38_combout ),
	.cout(\ram_rom_addr_reg[12]~39 ));
// synopsys translate_off
defparam \ram_rom_addr_reg[12]~38 .lut_mask = 16'hA50A;
defparam \ram_rom_addr_reg[12]~38 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X49_Y32_N28
cycloneive_lcell_comb \ram_rom_addr_reg[13]~40 (
	.dataa(gnd),
	.datab(ram_rom_addr_reg_13),
	.datac(gnd),
	.datad(gnd),
	.cin(\ram_rom_addr_reg[12]~39 ),
	.combout(\ram_rom_addr_reg[13]~40_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[13]~40 .lut_mask = 16'h3C3C;
defparam \ram_rom_addr_reg[13]~40 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N20
cycloneive_lcell_comb \process_0~3 (
	.dataa(node_ena_1),
	.datab(virtual_ir_scan_reg),
	.datac(ir_in[3]),
	.datad(state_4),
	.cin(gnd),
	.combout(\process_0~3_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~3 .lut_mask = 16'h2000;
defparam \process_0~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N30
cycloneive_lcell_comb \ram_rom_addr_reg[7]~42 (
	.dataa(\Equal1~1_combout ),
	.datab(\process_0~3_combout ),
	.datac(irf_reg_1_1),
	.datad(ram_rom_data_shift_cntr_reg[1]),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[7]~42_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~42 .lut_mask = 16'hCCEC;
defparam \ram_rom_addr_reg[7]~42 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N0
cycloneive_lcell_comb \ram_rom_addr_reg[7]~43 (
	.dataa(sdr),
	.datab(state_8),
	.datac(\ram_rom_addr_reg[7]~42_combout ),
	.datad(irf_reg_2_1),
	.cin(gnd),
	.combout(\ram_rom_addr_reg[7]~43_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_addr_reg[7]~43 .lut_mask = 16'hF8F0;
defparam \ram_rom_addr_reg[7]~43 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N14
cycloneive_lcell_comb \ram_rom_data_reg[1]~1 (
	.dataa(ram_block3a1),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a33),
	.cin(gnd),
	.combout(\ram_rom_data_reg[1]~1_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[1]~1 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[1]~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N8
cycloneive_lcell_comb \ram_rom_data_reg[2]~2 (
	.dataa(ram_block3a34),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a2),
	.cin(gnd),
	.combout(\ram_rom_data_reg[2]~2_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[2]~2 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[2]~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N22
cycloneive_lcell_comb \ram_rom_data_reg[3]~3 (
	.dataa(ram_block3a35),
	.datab(ram_block3a3),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[3]~3_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[3]~3 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[3]~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N24
cycloneive_lcell_comb \ram_rom_data_reg[4]~4 (
	.dataa(ram_block3a36),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a4),
	.cin(gnd),
	.combout(\ram_rom_data_reg[4]~4_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[4]~4 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[4]~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N24
cycloneive_lcell_comb \ram_rom_data_reg[5]~5 (
	.dataa(ram_block3a37),
	.datab(ram_block3a5),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[5]~5_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[5]~5 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[5]~5 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N18
cycloneive_lcell_comb \ram_rom_data_reg[6]~6 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a6),
	.datac(gnd),
	.datad(ram_block3a38),
	.cin(gnd),
	.combout(\ram_rom_data_reg[6]~6_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[6]~6 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[6]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N20
cycloneive_lcell_comb \ram_rom_data_reg[7]~7 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a39),
	.datac(gnd),
	.datad(ram_block3a7),
	.cin(gnd),
	.combout(\ram_rom_data_reg[7]~7_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[7]~7 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[7]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N30
cycloneive_lcell_comb \ram_rom_data_reg[8]~8 (
	.dataa(ram_block3a40),
	.datab(ram_block3a8),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[8]~8_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[8]~8 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[8]~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N16
cycloneive_lcell_comb \ram_rom_data_reg[9]~9 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a41),
	.datac(gnd),
	.datad(ram_block3a9),
	.cin(gnd),
	.combout(\ram_rom_data_reg[9]~9_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[9]~9 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[9]~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N10
cycloneive_lcell_comb \ram_rom_data_reg[10]~10 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a10),
	.datac(gnd),
	.datad(ram_block3a42),
	.cin(gnd),
	.combout(\ram_rom_data_reg[10]~10_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[10]~10 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[10]~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N28
cycloneive_lcell_comb \ram_rom_data_reg[11]~11 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a11),
	.datac(gnd),
	.datad(ram_block3a43),
	.cin(gnd),
	.combout(\ram_rom_data_reg[11]~11_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[11]~11 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[11]~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N26
cycloneive_lcell_comb \ram_rom_data_reg[12]~12 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a12),
	.datac(gnd),
	.datad(ram_block3a44),
	.cin(gnd),
	.combout(\ram_rom_data_reg[12]~12_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[12]~12 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[12]~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N8
cycloneive_lcell_comb \ram_rom_data_reg[13]~13 (
	.dataa(ram_block3a45),
	.datab(ram_block3a13),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[13]~13_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[13]~13 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[13]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X75_Y31_N14
cycloneive_lcell_comb \ram_rom_data_reg[14]~14 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a14),
	.datac(gnd),
	.datad(ram_block3a46),
	.cin(gnd),
	.combout(\ram_rom_data_reg[14]~14_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[14]~14 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[14]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N26
cycloneive_lcell_comb \ram_rom_data_reg[15]~15 (
	.dataa(ram_block3a47),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a15),
	.cin(gnd),
	.combout(\ram_rom_data_reg[15]~15_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[15]~15 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[15]~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N28
cycloneive_lcell_comb \ram_rom_data_reg[16]~16 (
	.dataa(ram_block3a48),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a16),
	.cin(gnd),
	.combout(\ram_rom_data_reg[16]~16_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[16]~16 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[16]~16 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N26
cycloneive_lcell_comb \ram_rom_data_reg[17]~17 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a49),
	.datac(gnd),
	.datad(ram_block3a17),
	.cin(gnd),
	.combout(\ram_rom_data_reg[17]~17_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[17]~17 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[17]~17 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N0
cycloneive_lcell_comb \ram_rom_data_reg[18]~18 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a50),
	.datac(gnd),
	.datad(ram_block3a18),
	.cin(gnd),
	.combout(\ram_rom_data_reg[18]~18_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[18]~18 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[18]~18 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N22
cycloneive_lcell_comb \ram_rom_data_reg[19]~19 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a19),
	.datac(gnd),
	.datad(ram_block3a51),
	.cin(gnd),
	.combout(\ram_rom_data_reg[19]~19_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[19]~19 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[19]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N8
cycloneive_lcell_comb \ram_rom_data_reg[20]~20 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a52),
	.datac(gnd),
	.datad(ram_block3a20),
	.cin(gnd),
	.combout(\ram_rom_data_reg[20]~20_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[20]~20 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[20]~20 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N18
cycloneive_lcell_comb \ram_rom_data_reg[21]~21 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a21),
	.datac(gnd),
	.datad(ram_block3a53),
	.cin(gnd),
	.combout(\ram_rom_data_reg[21]~21_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[21]~21 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[21]~21 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N4
cycloneive_lcell_comb \ram_rom_data_reg[22]~22 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a22),
	.datac(gnd),
	.datad(ram_block3a54),
	.cin(gnd),
	.combout(\ram_rom_data_reg[22]~22_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[22]~22 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[22]~22 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N30
cycloneive_lcell_comb \ram_rom_data_reg[23]~23 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a23),
	.datac(gnd),
	.datad(ram_block3a55),
	.cin(gnd),
	.combout(\ram_rom_data_reg[23]~23_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[23]~23 .lut_mask = 16'hEE44;
defparam \ram_rom_data_reg[23]~23 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N12
cycloneive_lcell_comb \ram_rom_data_reg[24]~24 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a56),
	.datac(gnd),
	.datad(ram_block3a24),
	.cin(gnd),
	.combout(\ram_rom_data_reg[24]~24_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[24]~24 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[24]~24 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N14
cycloneive_lcell_comb \ram_rom_data_reg[25]~25 (
	.dataa(address_reg_b_0),
	.datab(ram_block3a57),
	.datac(gnd),
	.datad(ram_block3a25),
	.cin(gnd),
	.combout(\ram_rom_data_reg[25]~25_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[25]~25 .lut_mask = 16'hDD88;
defparam \ram_rom_data_reg[25]~25 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X52_Y33_N20
cycloneive_lcell_comb \ram_rom_data_reg[26]~26 (
	.dataa(ram_block3a26),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a58),
	.cin(gnd),
	.combout(\ram_rom_data_reg[26]~26_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[26]~26 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[26]~26 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N12
cycloneive_lcell_comb \ram_rom_data_reg[27]~27 (
	.dataa(ram_block3a27),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a59),
	.cin(gnd),
	.combout(\ram_rom_data_reg[27]~27_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[27]~27 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[27]~27 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N18
cycloneive_lcell_comb \ram_rom_data_reg[28]~28 (
	.dataa(ram_block3a28),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a60),
	.cin(gnd),
	.combout(\ram_rom_data_reg[28]~28_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[28]~28 .lut_mask = 16'hEE22;
defparam \ram_rom_data_reg[28]~28 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N28
cycloneive_lcell_comb \ram_rom_data_reg[29]~29 (
	.dataa(ram_block3a61),
	.datab(ram_block3a29),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[29]~29_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[29]~29 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[29]~29 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N30
cycloneive_lcell_comb \ram_rom_data_reg[30]~30 (
	.dataa(ram_block3a62),
	.datab(address_reg_b_0),
	.datac(gnd),
	.datad(ram_block3a30),
	.cin(gnd),
	.combout(\ram_rom_data_reg[30]~30_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[30]~30 .lut_mask = 16'hBB88;
defparam \ram_rom_data_reg[30]~30 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X50_Y28_N16
cycloneive_lcell_comb \ram_rom_data_reg[31]~31 (
	.dataa(ram_block3a63),
	.datab(ram_block3a31),
	.datac(gnd),
	.datad(address_reg_b_0),
	.cin(gnd),
	.combout(\ram_rom_data_reg[31]~31_combout ),
	.cout());
// synopsys translate_off
defparam \ram_rom_data_reg[31]~31 .lut_mask = 16'hAACC;
defparam \ram_rom_data_reg[31]~31 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X47_Y32_N12
cycloneive_lcell_comb \process_0~0 (
	.dataa(ir_in[0]),
	.datab(gnd),
	.datac(irf_reg_4_1),
	.datad(gnd),
	.cin(gnd),
	.combout(\process_0~0_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~0 .lut_mask = 16'hFAFA;
defparam \process_0~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N26
cycloneive_lcell_comb \process_0~1 (
	.dataa(virtual_ir_scan_reg),
	.datab(ir_in[3]),
	.datac(state_5),
	.datad(node_ena_1),
	.cin(gnd),
	.combout(\process_0~1_combout ),
	.cout());
// synopsys translate_off
defparam \process_0~1 .lut_mask = 16'h4000;
defparam \process_0~1 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N2
cycloneive_lcell_comb \ir_loaded_address_reg[1]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_1),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[1]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[1]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[1]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N24
cycloneive_lcell_comb \ir_loaded_address_reg[2]~feeder (
	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(ram_rom_addr_reg_2),
	.cin(gnd),
	.combout(\ir_loaded_address_reg[2]~feeder_combout ),
	.cout());
// synopsys translate_off
defparam \ir_loaded_address_reg[2]~feeder .lut_mask = 16'hFF00;
defparam \ir_loaded_address_reg[2]~feeder .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N28
cycloneive_lcell_comb \bypass_reg_out~0 (
	.dataa(altera_internal_jtag),
	.datab(gnd),
	.datac(\bypass_reg_out~q ),
	.datad(node_ena_1),
	.cin(gnd),
	.combout(\bypass_reg_out~0_combout ),
	.cout());
// synopsys translate_off
defparam \bypass_reg_out~0 .lut_mask = 16'hAAF0;
defparam \bypass_reg_out~0 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X46_Y32_N29
dffeas bypass_reg_out(
	.clk(raw_tck),
	.d(\bypass_reg_out~0_combout ),
	.asdata(vcc),
	.clrn(!clr),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(\bypass_reg_out~q ),
	.prn(vcc));
// synopsys translate_off
defparam bypass_reg_out.is_wysiwyg = "true";
defparam bypass_reg_out.power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X46_Y32_N14
cycloneive_lcell_comb \tdo~0 (
	.dataa(irf_reg_1_1),
	.datab(irf_reg_2_1),
	.datac(ram_rom_data_reg_0),
	.datad(\bypass_reg_out~q ),
	.cin(gnd),
	.combout(\tdo~0_combout ),
	.cout());
// synopsys translate_off
defparam \tdo~0 .lut_mask = 16'hF1E0;
defparam \tdo~0 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule

module sld_rom_sr (
	WORD_SR_0,
	sdr,
	altera_internal_jtag,
	state_4,
	virtual_ir_scan_reg,
	state_3,
	state_8,
	TCK,
	devpor,
	devclrn,
	devoe);
output 	WORD_SR_0;
input 	sdr;
input 	altera_internal_jtag;
input 	state_4;
input 	virtual_ir_scan_reg;
input 	state_3;
input 	state_8;
input 	TCK;

// Design Ports Information

input 	devpor;
input 	devclrn;
input 	devoe;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

wire \WORD_SR~7_combout ;
wire \WORD_SR~8_combout ;
wire \WORD_SR~10_combout ;
wire \WORD_SR~11_combout ;
wire \WORD_SR~13_combout ;
wire \word_counter[0]~7_combout ;
wire \word_counter[0]~8 ;
wire \word_counter[1]~9_combout ;
wire \clear_signal~combout ;
wire \word_counter[0]~14_combout ;
wire \word_counter[1]~10 ;
wire \word_counter[2]~11_combout ;
wire \word_counter[2]~12 ;
wire \word_counter[3]~15_combout ;
wire \word_counter[3]~16 ;
wire \word_counter[4]~17_combout ;
wire \word_counter[0]~13_combout ;
wire \word_counter[0]~19_combout ;
wire \WORD_SR~14_combout ;
wire \WORD_SR~15_combout ;
wire \WORD_SR[3]~6_combout ;
wire \WORD_SR~12_combout ;
wire \WORD_SR~9_combout ;
wire \WORD_SR~3_combout ;
wire \WORD_SR~2_combout ;
wire \WORD_SR~4_combout ;
wire \WORD_SR~5_combout ;
wire [4:0] word_counter;
wire [3:0] WORD_SR;


// Location: LCCOMB_X43_Y32_N22
cycloneive_lcell_comb \WORD_SR~7 (
	.dataa(word_counter[1]),
	.datab(state_4),
	.datac(word_counter[0]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~7_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~7 .lut_mask = 16'h0203;
defparam \WORD_SR~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N12
cycloneive_lcell_comb \WORD_SR~8 (
	.dataa(\WORD_SR~7_combout ),
	.datab(word_counter[2]),
	.datac(word_counter[3]),
	.datad(gnd),
	.cin(gnd),
	.combout(\WORD_SR~8_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~8 .lut_mask = 16'h0202;
defparam \WORD_SR~8 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N26
cycloneive_lcell_comb \WORD_SR~10 (
	.dataa(word_counter[2]),
	.datab(word_counter[0]),
	.datac(word_counter[4]),
	.datad(word_counter[1]),
	.cin(gnd),
	.combout(\WORD_SR~10_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~10 .lut_mask = 16'hD8F2;
defparam \WORD_SR~10 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N12
cycloneive_lcell_comb \WORD_SR~11 (
	.dataa(gnd),
	.datab(word_counter[0]),
	.datac(\WORD_SR~10_combout ),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~11_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~11 .lut_mask = 16'hC3C0;
defparam \WORD_SR~11 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N30
cycloneive_lcell_comb \WORD_SR~13 (
	.dataa(word_counter[1]),
	.datab(word_counter[2]),
	.datac(word_counter[3]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~13_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~13 .lut_mask = 16'h0080;
defparam \WORD_SR~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N29
dffeas \WORD_SR[0] (
	.clk(TCK),
	.d(\WORD_SR~5_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR_0),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[0] .is_wysiwyg = "true";
defparam \WORD_SR[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N0
cycloneive_lcell_comb \word_counter[0]~7 (
	.dataa(gnd),
	.datab(word_counter[0]),
	.datac(gnd),
	.datad(vcc),
	.cin(gnd),
	.combout(\word_counter[0]~7_combout ),
	.cout(\word_counter[0]~8 ));
// synopsys translate_off
defparam \word_counter[0]~7 .lut_mask = 16'h33CC;
defparam \word_counter[0]~7 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N2
cycloneive_lcell_comb \word_counter[1]~9 (
	.dataa(gnd),
	.datab(word_counter[1]),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[0]~8 ),
	.combout(\word_counter[1]~9_combout ),
	.cout(\word_counter[1]~10 ));
// synopsys translate_off
defparam \word_counter[1]~9 .lut_mask = 16'h3C3F;
defparam \word_counter[1]~9 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N8
cycloneive_lcell_comb clear_signal(
	.dataa(gnd),
	.datab(gnd),
	.datac(state_8),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\clear_signal~combout ),
	.cout());
// synopsys translate_off
defparam clear_signal.lut_mask = 16'hF000;
defparam clear_signal.sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N18
cycloneive_lcell_comb \word_counter[0]~14 (
	.dataa(sdr),
	.datab(\clear_signal~combout ),
	.datac(state_3),
	.datad(state_4),
	.cin(gnd),
	.combout(\word_counter[0]~14_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[0]~14 .lut_mask = 16'hCCEC;
defparam \word_counter[0]~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y32_N3
dffeas \word_counter[1] (
	.clk(TCK),
	.d(\word_counter[1]~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[1]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[1] .is_wysiwyg = "true";
defparam \word_counter[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N4
cycloneive_lcell_comb \word_counter[2]~11 (
	.dataa(word_counter[2]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[1]~10 ),
	.combout(\word_counter[2]~11_combout ),
	.cout(\word_counter[2]~12 ));
// synopsys translate_off
defparam \word_counter[2]~11 .lut_mask = 16'hA50A;
defparam \word_counter[2]~11 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X42_Y32_N5
dffeas \word_counter[2] (
	.clk(TCK),
	.d(\word_counter[2]~11_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[2]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[2] .is_wysiwyg = "true";
defparam \word_counter[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N6
cycloneive_lcell_comb \word_counter[3]~15 (
	.dataa(word_counter[3]),
	.datab(gnd),
	.datac(gnd),
	.datad(vcc),
	.cin(\word_counter[2]~12 ),
	.combout(\word_counter[3]~15_combout ),
	.cout(\word_counter[3]~16 ));
// synopsys translate_off
defparam \word_counter[3]~15 .lut_mask = 16'h5A5F;
defparam \word_counter[3]~15 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X42_Y32_N7
dffeas \word_counter[3] (
	.clk(TCK),
	.d(\word_counter[3]~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[3]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[3] .is_wysiwyg = "true";
defparam \word_counter[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X42_Y32_N8
cycloneive_lcell_comb \word_counter[4]~17 (
	.dataa(gnd),
	.datab(word_counter[4]),
	.datac(gnd),
	.datad(gnd),
	.cin(\word_counter[3]~16 ),
	.combout(\word_counter[4]~17_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[4]~17 .lut_mask = 16'hC3C3;
defparam \word_counter[4]~17 .sum_lutc_input = "cin";
// synopsys translate_on

// Location: FF_X42_Y32_N9
dffeas \word_counter[4] (
	.clk(TCK),
	.d(\word_counter[4]~17_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[4]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[4] .is_wysiwyg = "true";
defparam \word_counter[4] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N24
cycloneive_lcell_comb \word_counter[0]~13 (
	.dataa(word_counter[1]),
	.datab(word_counter[2]),
	.datac(word_counter[3]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\word_counter[0]~13_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[0]~13 .lut_mask = 16'hFBFF;
defparam \word_counter[0]~13 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N26
cycloneive_lcell_comb \word_counter[0]~19 (
	.dataa(word_counter[0]),
	.datab(\word_counter[0]~13_combout ),
	.datac(state_8),
	.datad(virtual_ir_scan_reg),
	.cin(gnd),
	.combout(\word_counter[0]~19_combout ),
	.cout());
// synopsys translate_off
defparam \word_counter[0]~19 .lut_mask = 16'hF111;
defparam \word_counter[0]~19 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X42_Y32_N1
dffeas \word_counter[0] (
	.clk(TCK),
	.d(\word_counter[0]~7_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(\word_counter[0]~19_combout ),
	.sload(gnd),
	.ena(\word_counter[0]~14_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(word_counter[0]),
	.prn(vcc));
// synopsys translate_off
defparam \word_counter[0] .is_wysiwyg = "true";
defparam \word_counter[0] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N20
cycloneive_lcell_comb \WORD_SR~14 (
	.dataa(\WORD_SR~13_combout ),
	.datab(altera_internal_jtag),
	.datac(word_counter[0]),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~14_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~14 .lut_mask = 16'hCC0A;
defparam \WORD_SR~14 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N0
cycloneive_lcell_comb \WORD_SR~15 (
	.dataa(virtual_ir_scan_reg),
	.datab(gnd),
	.datac(state_8),
	.datad(\WORD_SR~14_combout ),
	.cin(gnd),
	.combout(\WORD_SR~15_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~15 .lut_mask = 16'h5F00;
defparam \WORD_SR~15 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N16
cycloneive_lcell_comb \WORD_SR[3]~6 (
	.dataa(sdr),
	.datab(\clear_signal~combout ),
	.datac(state_3),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR[3]~6_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR[3]~6 .lut_mask = 16'hEEEC;
defparam \WORD_SR[3]~6 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N1
dffeas \WORD_SR[3] (
	.clk(TCK),
	.d(\WORD_SR~15_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[3]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[3] .is_wysiwyg = "true";
defparam \WORD_SR[3] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N2
cycloneive_lcell_comb \WORD_SR~12 (
	.dataa(\WORD_SR~11_combout ),
	.datab(WORD_SR[3]),
	.datac(\clear_signal~combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~12_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~12 .lut_mask = 16'h0C0A;
defparam \WORD_SR~12 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N3
dffeas \WORD_SR[2] (
	.clk(TCK),
	.d(\WORD_SR~12_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[2]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[2] .is_wysiwyg = "true";
defparam \WORD_SR[2] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N10
cycloneive_lcell_comb \WORD_SR~9 (
	.dataa(\WORD_SR~8_combout ),
	.datab(WORD_SR[2]),
	.datac(\clear_signal~combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~9_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~9 .lut_mask = 16'h0E0A;
defparam \WORD_SR~9 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: FF_X43_Y32_N11
dffeas \WORD_SR[1] (
	.clk(TCK),
	.d(\WORD_SR~9_combout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(\WORD_SR[3]~6_combout ),
	.devclrn(devclrn),
	.devpor(devpor),
	.q(WORD_SR[1]),
	.prn(vcc));
// synopsys translate_off
defparam \WORD_SR[1] .is_wysiwyg = "true";
defparam \WORD_SR[1] .power_up = "low";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N4
cycloneive_lcell_comb \WORD_SR~3 (
	.dataa(word_counter[1]),
	.datab(word_counter[2]),
	.datac(word_counter[0]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~3_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~3 .lut_mask = 16'hAB08;
defparam \WORD_SR~3 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N6
cycloneive_lcell_comb \WORD_SR~2 (
	.dataa(word_counter[1]),
	.datab(word_counter[2]),
	.datac(word_counter[3]),
	.datad(word_counter[4]),
	.cin(gnd),
	.combout(\WORD_SR~2_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~2 .lut_mask = 16'h01C1;
defparam \WORD_SR~2 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N14
cycloneive_lcell_comb \WORD_SR~4 (
	.dataa(gnd),
	.datab(\WORD_SR~3_combout ),
	.datac(word_counter[0]),
	.datad(\WORD_SR~2_combout ),
	.cin(gnd),
	.combout(\WORD_SR~4_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~4 .lut_mask = 16'hCCC0;
defparam \WORD_SR~4 .sum_lutc_input = "datac";
// synopsys translate_on

// Location: LCCOMB_X43_Y32_N28
cycloneive_lcell_comb \WORD_SR~5 (
	.dataa(WORD_SR[1]),
	.datab(\WORD_SR~4_combout ),
	.datac(\clear_signal~combout ),
	.datad(state_4),
	.cin(gnd),
	.combout(\WORD_SR~5_combout ),
	.cout());
// synopsys translate_off
defparam \WORD_SR~5 .lut_mask = 16'h0A0C;
defparam \WORD_SR~5 .sum_lutc_input = "datac";
// synopsys translate_on

endmodule
